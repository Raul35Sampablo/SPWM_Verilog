module mem2(

	input clk,									//señal de reloj
	//input reset_mem2,							
	input  [14:0] selector2,				//seleccion de ubicacion de memoria
	output reg[9:0] output_data_2 		//salida de nuestra onda senoidal en señal

);
reg [9:0] mem2 [0:15359];

initial begin
mem2[0] = 10'b0000000000;
mem2[1] = 10'b0000000000;
mem2[2] = 10'b0000000000;
mem2[3] = 10'b0000000000;
mem2[4] = 10'b0000000000;
mem2[5] = 10'b0000000000;
mem2[6] = 10'b0000000000;
mem2[7] = 10'b0000000000;
mem2[8] = 10'b0000000000;
mem2[9] = 10'b0000000000;
mem2[10] = 10'b0000000000;
mem2[11] = 10'b0000000000;
mem2[12] = 10'b0000000000;
mem2[13] = 10'b0000000000;
mem2[14] = 10'b0000000000;
mem2[15] = 10'b0000000000;
mem2[16] = 10'b0000000000;
mem2[17] = 10'b0000000000;
mem2[18] = 10'b0000000000;
mem2[19] = 10'b0000000000;
mem2[20] = 10'b0000000000;
mem2[21] = 10'b0000000000;
mem2[22] = 10'b0000000000;
mem2[23] = 10'b0000000000;
mem2[24] = 10'b0000000000;
mem2[25] = 10'b0000000000;
mem2[26] = 10'b0000000000;
mem2[27] = 10'b0000000000;
mem2[28] = 10'b0000000000;
mem2[29] = 10'b0000000000;
mem2[30] = 10'b0000000000;
mem2[31] = 10'b0000000000;
mem2[32] = 10'b0000000000;
mem2[33] = 10'b0000000000;
mem2[34] = 10'b0000000000;
mem2[35] = 10'b0000000000;
mem2[36] = 10'b0000000000;
mem2[37] = 10'b0000000000;
mem2[38] = 10'b0000000000;
mem2[39] = 10'b0000000000;
mem2[40] = 10'b0000000000;
mem2[41] = 10'b0000000000;
mem2[42] = 10'b0000000000;
mem2[43] = 10'b0000000000;
mem2[44] = 10'b0000000000;
mem2[45] = 10'b0000000000;
mem2[46] = 10'b0000000000;
mem2[47] = 10'b0000000000;
mem2[48] = 10'b0000000000;
mem2[49] = 10'b0000000000;
mem2[50] = 10'b0000000000;
mem2[51] = 10'b0000000000;
mem2[52] = 10'b0000000000;
mem2[53] = 10'b0000000000;
mem2[54] = 10'b0000000000;
mem2[55] = 10'b0000000000;
mem2[56] = 10'b0000000000;
mem2[57] = 10'b0000000000;
mem2[58] = 10'b0000000000;
mem2[59] = 10'b0000000000;
mem2[60] = 10'b0000000000;
mem2[61] = 10'b0000000000;
mem2[62] = 10'b0000000000;
mem2[63] = 10'b0000000000;
mem2[64] = 10'b0000000000;
mem2[65] = 10'b0000000000;
mem2[66] = 10'b0000000000;
mem2[67] = 10'b0000000000;
mem2[68] = 10'b0000000000;
mem2[69] = 10'b0000000000;
mem2[70] = 10'b0000000000;
mem2[71] = 10'b0000000000;
mem2[72] = 10'b0000000000;
mem2[73] = 10'b0000000000;
mem2[74] = 10'b0000000000;
mem2[75] = 10'b0000000000;
mem2[76] = 10'b0000000000;
mem2[77] = 10'b0000000000;
mem2[78] = 10'b0000000000;
mem2[79] = 10'b0000000000;
mem2[80] = 10'b0000000000;
mem2[81] = 10'b0000000000;
mem2[82] = 10'b0000000000;
mem2[83] = 10'b0000000000;
mem2[84] = 10'b0000000000;
mem2[85] = 10'b0000000000;
mem2[86] = 10'b0000000000;
mem2[87] = 10'b0000000000;
mem2[88] = 10'b0000000000;
mem2[89] = 10'b0000000000;
mem2[90] = 10'b0000000000;
mem2[91] = 10'b0000000000;
mem2[92] = 10'b0000000000;
mem2[93] = 10'b0000000000;
mem2[94] = 10'b0000000000;
mem2[95] = 10'b0000000000;
mem2[96] = 10'b0000000000;
mem2[97] = 10'b0000000000;
mem2[98] = 10'b0000000000;
mem2[99] = 10'b0000000000;
mem2[100] = 10'b0000000000;
mem2[101] = 10'b0000000000;
mem2[102] = 10'b0000000000;
mem2[103] = 10'b0000000000;
mem2[104] = 10'b0000000000;
mem2[105] = 10'b0000000000;
mem2[106] = 10'b0000000000;
mem2[107] = 10'b0000000000;
mem2[108] = 10'b0000000000;
mem2[109] = 10'b0000000000;
mem2[110] = 10'b0000000000;
mem2[111] = 10'b0000000000;
mem2[112] = 10'b0000000000;
mem2[113] = 10'b0000000000;
mem2[114] = 10'b0000000000;
mem2[115] = 10'b0000000000;
mem2[116] = 10'b0000000000;
mem2[117] = 10'b0000000000;
mem2[118] = 10'b0000000000;
mem2[119] = 10'b0000000000;
mem2[120] = 10'b0000000000;
mem2[121] = 10'b0000000000;
mem2[122] = 10'b0000000000;
mem2[123] = 10'b0000000000;
mem2[124] = 10'b0000000000;
mem2[125] = 10'b0000000000;
mem2[126] = 10'b0000000000;
mem2[127] = 10'b0000000000;
mem2[128] = 10'b0000000000;
mem2[129] = 10'b0000000000;
mem2[130] = 10'b0000000000;
mem2[131] = 10'b0000000000;
mem2[132] = 10'b0000000000;
mem2[133] = 10'b0000000000;
mem2[134] = 10'b0000000000;
mem2[135] = 10'b0000000000;
mem2[136] = 10'b0000000000;
mem2[137] = 10'b0000000000;
mem2[138] = 10'b0000000000;
mem2[139] = 10'b0000000000;
mem2[140] = 10'b0000000000;
mem2[141] = 10'b0000000000;
mem2[142] = 10'b0000000000;
mem2[143] = 10'b0000000000;
mem2[144] = 10'b0000000000;
mem2[145] = 10'b0000000000;
mem2[146] = 10'b0000000000;
mem2[147] = 10'b0000000000;
mem2[148] = 10'b0000000000;
mem2[149] = 10'b0000000000;
mem2[150] = 10'b0000000000;
mem2[151] = 10'b0000000000;
mem2[152] = 10'b0000000000;
mem2[153] = 10'b0000000000;
mem2[154] = 10'b0000000000;
mem2[155] = 10'b0000000000;
mem2[156] = 10'b0000000000;
mem2[157] = 10'b0000000000;
mem2[158] = 10'b0000000000;
mem2[159] = 10'b0000000000;
mem2[160] = 10'b0000000000;
mem2[161] = 10'b0000000000;
mem2[162] = 10'b0000000000;
mem2[163] = 10'b0000000000;
mem2[164] = 10'b0000000000;
mem2[165] = 10'b0000000000;
mem2[166] = 10'b0000000000;
mem2[167] = 10'b0000000000;
mem2[168] = 10'b0000000000;
mem2[169] = 10'b0000000000;
mem2[170] = 10'b0000000000;
mem2[171] = 10'b0000000000;
mem2[172] = 10'b0000000000;
mem2[173] = 10'b0000000000;
mem2[174] = 10'b0000000000;
mem2[175] = 10'b0000000000;
mem2[176] = 10'b0000000000;
mem2[177] = 10'b0000000000;
mem2[178] = 10'b0000000000;
mem2[179] = 10'b0000000000;
mem2[180] = 10'b0000000000;
mem2[181] = 10'b0000000000;
mem2[182] = 10'b0000000000;
mem2[183] = 10'b0000000000;
mem2[184] = 10'b0000000000;
mem2[185] = 10'b0000000000;
mem2[186] = 10'b0000000000;
mem2[187] = 10'b0000000000;
mem2[188] = 10'b0000000000;
mem2[189] = 10'b0000000000;
mem2[190] = 10'b0000000000;
mem2[191] = 10'b0000000000;
mem2[192] = 10'b0000000000;
mem2[193] = 10'b0000000000;
mem2[194] = 10'b0000000000;
mem2[195] = 10'b0000000000;
mem2[196] = 10'b0000000000;
mem2[197] = 10'b0000000000;
mem2[198] = 10'b0000000000;
mem2[199] = 10'b0000000000;
mem2[200] = 10'b0000000000;
mem2[201] = 10'b0000000000;
mem2[202] = 10'b0000000000;
mem2[203] = 10'b0000000000;
mem2[204] = 10'b0000000000;
mem2[205] = 10'b0000000000;
mem2[206] = 10'b0000000000;
mem2[207] = 10'b0000000000;
mem2[208] = 10'b0000000000;
mem2[209] = 10'b0000000000;
mem2[210] = 10'b0000000000;
mem2[211] = 10'b0000000000;
mem2[212] = 10'b0000000000;
mem2[213] = 10'b0000000000;
mem2[214] = 10'b0000000000;
mem2[215] = 10'b0000000000;
mem2[216] = 10'b0000000000;
mem2[217] = 10'b0000000000;
mem2[218] = 10'b0000000000;
mem2[219] = 10'b0000000000;
mem2[220] = 10'b0000000000;
mem2[221] = 10'b0000000000;
mem2[222] = 10'b0000000000;
mem2[223] = 10'b0000000000;
mem2[224] = 10'b0000000000;
mem2[225] = 10'b0000000000;
mem2[226] = 10'b0000000000;
mem2[227] = 10'b0000000000;
mem2[228] = 10'b0000000000;
mem2[229] = 10'b0000000000;
mem2[230] = 10'b0000000000;
mem2[231] = 10'b0000000000;
mem2[232] = 10'b0000000000;
mem2[233] = 10'b0000000000;
mem2[234] = 10'b0000000000;
mem2[235] = 10'b0000000000;
mem2[236] = 10'b0000000000;
mem2[237] = 10'b0000000000;
mem2[238] = 10'b0000000000;
mem2[239] = 10'b0000000000;
mem2[240] = 10'b0000000000;
mem2[241] = 10'b0000000000;
mem2[242] = 10'b0000000000;
mem2[243] = 10'b0000000000;
mem2[244] = 10'b0000000000;
mem2[245] = 10'b0000000000;
mem2[246] = 10'b0000000000;
mem2[247] = 10'b0000000000;
mem2[248] = 10'b0000000000;
mem2[249] = 10'b0000000000;
mem2[250] = 10'b0000000000;
mem2[251] = 10'b0000000000;
mem2[252] = 10'b0000000000;
mem2[253] = 10'b0000000000;
mem2[254] = 10'b0000000000;
mem2[255] = 10'b0000000000;
mem2[256] = 10'b0000000000;
mem2[257] = 10'b0000000000;
mem2[258] = 10'b0000000000;
mem2[259] = 10'b0000000000;
mem2[260] = 10'b0000000000;
mem2[261] = 10'b0000000000;
mem2[262] = 10'b0000000000;
mem2[263] = 10'b0000000000;
mem2[264] = 10'b0000000000;
mem2[265] = 10'b0000000000;
mem2[266] = 10'b0000000000;
mem2[267] = 10'b0000000000;
mem2[268] = 10'b0000000000;
mem2[269] = 10'b0000000000;
mem2[270] = 10'b0000000000;
mem2[271] = 10'b0000000000;
mem2[272] = 10'b0000000000;
mem2[273] = 10'b0000000000;
mem2[274] = 10'b0000000000;
mem2[275] = 10'b0000000000;
mem2[276] = 10'b0000000000;
mem2[277] = 10'b0000000000;
mem2[278] = 10'b0000000000;
mem2[279] = 10'b0000000000;
mem2[280] = 10'b0000000000;
mem2[281] = 10'b0000000000;
mem2[282] = 10'b0000000000;
mem2[283] = 10'b0000000000;
mem2[284] = 10'b0000000000;
mem2[285] = 10'b0000000000;
mem2[286] = 10'b0000000000;
mem2[287] = 10'b0000000000;
mem2[288] = 10'b0000000000;
mem2[289] = 10'b0000000000;
mem2[290] = 10'b0000000000;
mem2[291] = 10'b0000000000;
mem2[292] = 10'b0000000000;
mem2[293] = 10'b0000000000;
mem2[294] = 10'b0000000000;
mem2[295] = 10'b0000000000;
mem2[296] = 10'b0000000000;
mem2[297] = 10'b0000000000;
mem2[298] = 10'b0000000000;
mem2[299] = 10'b0000000000;
mem2[300] = 10'b0000000000;
mem2[301] = 10'b0000000000;
mem2[302] = 10'b0000000000;
mem2[303] = 10'b0000000000;
mem2[304] = 10'b0000000000;
mem2[305] = 10'b0000000000;
mem2[306] = 10'b0000000001;
mem2[307] = 10'b0000000001;
mem2[308] = 10'b0000000001;
mem2[309] = 10'b0000000001;
mem2[310] = 10'b0000000001;
mem2[311] = 10'b0000000001;
mem2[312] = 10'b0000000001;
mem2[313] = 10'b0000000001;
mem2[314] = 10'b0000000001;
mem2[315] = 10'b0000000001;
mem2[316] = 10'b0000000001;
mem2[317] = 10'b0000000001;
mem2[318] = 10'b0000000001;
mem2[319] = 10'b0000000001;
mem2[320] = 10'b0000000001;
mem2[321] = 10'b0000000001;
mem2[322] = 10'b0000000001;
mem2[323] = 10'b0000000001;
mem2[324] = 10'b0000000001;
mem2[325] = 10'b0000000001;
mem2[326] = 10'b0000000001;
mem2[327] = 10'b0000000001;
mem2[328] = 10'b0000000001;
mem2[329] = 10'b0000000001;
mem2[330] = 10'b0000000001;
mem2[331] = 10'b0000000001;
mem2[332] = 10'b0000000001;
mem2[333] = 10'b0000000001;
mem2[334] = 10'b0000000001;
mem2[335] = 10'b0000000001;
mem2[336] = 10'b0000000001;
mem2[337] = 10'b0000000001;
mem2[338] = 10'b0000000001;
mem2[339] = 10'b0000000001;
mem2[340] = 10'b0000000001;
mem2[341] = 10'b0000000001;
mem2[342] = 10'b0000000001;
mem2[343] = 10'b0000000001;
mem2[344] = 10'b0000000001;
mem2[345] = 10'b0000000001;
mem2[346] = 10'b0000000001;
mem2[347] = 10'b0000000001;
mem2[348] = 10'b0000000001;
mem2[349] = 10'b0000000001;
mem2[350] = 10'b0000000001;
mem2[351] = 10'b0000000001;
mem2[352] = 10'b0000000001;
mem2[353] = 10'b0000000001;
mem2[354] = 10'b0000000001;
mem2[355] = 10'b0000000001;
mem2[356] = 10'b0000000001;
mem2[357] = 10'b0000000001;
mem2[358] = 10'b0000000001;
mem2[359] = 10'b0000000001;
mem2[360] = 10'b0000000001;
mem2[361] = 10'b0000000001;
mem2[362] = 10'b0000000001;
mem2[363] = 10'b0000000001;
mem2[364] = 10'b0000000001;
mem2[365] = 10'b0000000001;
mem2[366] = 10'b0000000001;
mem2[367] = 10'b0000000001;
mem2[368] = 10'b0000000001;
mem2[369] = 10'b0000000001;
mem2[370] = 10'b0000000001;
mem2[371] = 10'b0000000001;
mem2[372] = 10'b0000000001;
mem2[373] = 10'b0000000001;
mem2[374] = 10'b0000000001;
mem2[375] = 10'b0000000001;
mem2[376] = 10'b0000000001;
mem2[377] = 10'b0000000001;
mem2[378] = 10'b0000000001;
mem2[379] = 10'b0000000001;
mem2[380] = 10'b0000000001;
mem2[381] = 10'b0000000001;
mem2[382] = 10'b0000000001;
mem2[383] = 10'b0000000001;
mem2[384] = 10'b0000000001;
mem2[385] = 10'b0000000001;
mem2[386] = 10'b0000000001;
mem2[387] = 10'b0000000001;
mem2[388] = 10'b0000000001;
mem2[389] = 10'b0000000001;
mem2[390] = 10'b0000000001;
mem2[391] = 10'b0000000001;
mem2[392] = 10'b0000000001;
mem2[393] = 10'b0000000001;
mem2[394] = 10'b0000000001;
mem2[395] = 10'b0000000001;
mem2[396] = 10'b0000000001;
mem2[397] = 10'b0000000001;
mem2[398] = 10'b0000000001;
mem2[399] = 10'b0000000001;
mem2[400] = 10'b0000000001;
mem2[401] = 10'b0000000001;
mem2[402] = 10'b0000000001;
mem2[403] = 10'b0000000001;
mem2[404] = 10'b0000000001;
mem2[405] = 10'b0000000001;
mem2[406] = 10'b0000000001;
mem2[407] = 10'b0000000001;
mem2[408] = 10'b0000000001;
mem2[409] = 10'b0000000001;
mem2[410] = 10'b0000000001;
mem2[411] = 10'b0000000001;
mem2[412] = 10'b0000000001;
mem2[413] = 10'b0000000001;
mem2[414] = 10'b0000000001;
mem2[415] = 10'b0000000001;
mem2[416] = 10'b0000000001;
mem2[417] = 10'b0000000001;
mem2[418] = 10'b0000000001;
mem2[419] = 10'b0000000001;
mem2[420] = 10'b0000000001;
mem2[421] = 10'b0000000001;
mem2[422] = 10'b0000000001;
mem2[423] = 10'b0000000001;
mem2[424] = 10'b0000000001;
mem2[425] = 10'b0000000001;
mem2[426] = 10'b0000000001;
mem2[427] = 10'b0000000001;
mem2[428] = 10'b0000000001;
mem2[429] = 10'b0000000001;
mem2[430] = 10'b0000000001;
mem2[431] = 10'b0000000001;
mem2[432] = 10'b0000000001;
mem2[433] = 10'b0000000010;
mem2[434] = 10'b0000000010;
mem2[435] = 10'b0000000010;
mem2[436] = 10'b0000000010;
mem2[437] = 10'b0000000010;
mem2[438] = 10'b0000000010;
mem2[439] = 10'b0000000010;
mem2[440] = 10'b0000000010;
mem2[441] = 10'b0000000010;
mem2[442] = 10'b0000000010;
mem2[443] = 10'b0000000010;
mem2[444] = 10'b0000000010;
mem2[445] = 10'b0000000010;
mem2[446] = 10'b0000000010;
mem2[447] = 10'b0000000010;
mem2[448] = 10'b0000000010;
mem2[449] = 10'b0000000010;
mem2[450] = 10'b0000000010;
mem2[451] = 10'b0000000010;
mem2[452] = 10'b0000000010;
mem2[453] = 10'b0000000010;
mem2[454] = 10'b0000000010;
mem2[455] = 10'b0000000010;
mem2[456] = 10'b0000000010;
mem2[457] = 10'b0000000010;
mem2[458] = 10'b0000000010;
mem2[459] = 10'b0000000010;
mem2[460] = 10'b0000000010;
mem2[461] = 10'b0000000010;
mem2[462] = 10'b0000000010;
mem2[463] = 10'b0000000010;
mem2[464] = 10'b0000000010;
mem2[465] = 10'b0000000010;
mem2[466] = 10'b0000000010;
mem2[467] = 10'b0000000010;
mem2[468] = 10'b0000000010;
mem2[469] = 10'b0000000010;
mem2[470] = 10'b0000000010;
mem2[471] = 10'b0000000010;
mem2[472] = 10'b0000000010;
mem2[473] = 10'b0000000010;
mem2[474] = 10'b0000000010;
mem2[475] = 10'b0000000010;
mem2[476] = 10'b0000000010;
mem2[477] = 10'b0000000010;
mem2[478] = 10'b0000000010;
mem2[479] = 10'b0000000010;
mem2[480] = 10'b0000000010;
mem2[481] = 10'b0000000010;
mem2[482] = 10'b0000000010;
mem2[483] = 10'b0000000010;
mem2[484] = 10'b0000000010;
mem2[485] = 10'b0000000010;
mem2[486] = 10'b0000000010;
mem2[487] = 10'b0000000010;
mem2[488] = 10'b0000000010;
mem2[489] = 10'b0000000010;
mem2[490] = 10'b0000000010;
mem2[491] = 10'b0000000010;
mem2[492] = 10'b0000000010;
mem2[493] = 10'b0000000010;
mem2[494] = 10'b0000000010;
mem2[495] = 10'b0000000010;
mem2[496] = 10'b0000000010;
mem2[497] = 10'b0000000010;
mem2[498] = 10'b0000000010;
mem2[499] = 10'b0000000010;
mem2[500] = 10'b0000000010;
mem2[501] = 10'b0000000010;
mem2[502] = 10'b0000000010;
mem2[503] = 10'b0000000010;
mem2[504] = 10'b0000000010;
mem2[505] = 10'b0000000010;
mem2[506] = 10'b0000000010;
mem2[507] = 10'b0000000010;
mem2[508] = 10'b0000000010;
mem2[509] = 10'b0000000010;
mem2[510] = 10'b0000000010;
mem2[511] = 10'b0000000010;
mem2[512] = 10'b0000000010;
mem2[513] = 10'b0000000010;
mem2[514] = 10'b0000000010;
mem2[515] = 10'b0000000010;
mem2[516] = 10'b0000000010;
mem2[517] = 10'b0000000010;
mem2[518] = 10'b0000000010;
mem2[519] = 10'b0000000010;
mem2[520] = 10'b0000000010;
mem2[521] = 10'b0000000010;
mem2[522] = 10'b0000000010;
mem2[523] = 10'b0000000010;
mem2[524] = 10'b0000000010;
mem2[525] = 10'b0000000010;
mem2[526] = 10'b0000000010;
mem2[527] = 10'b0000000010;
mem2[528] = 10'b0000000010;
mem2[529] = 10'b0000000010;
mem2[530] = 10'b0000000011;
mem2[531] = 10'b0000000011;
mem2[532] = 10'b0000000011;
mem2[533] = 10'b0000000011;
mem2[534] = 10'b0000000011;
mem2[535] = 10'b0000000011;
mem2[536] = 10'b0000000011;
mem2[537] = 10'b0000000011;
mem2[538] = 10'b0000000011;
mem2[539] = 10'b0000000011;
mem2[540] = 10'b0000000011;
mem2[541] = 10'b0000000011;
mem2[542] = 10'b0000000011;
mem2[543] = 10'b0000000011;
mem2[544] = 10'b0000000011;
mem2[545] = 10'b0000000011;
mem2[546] = 10'b0000000011;
mem2[547] = 10'b0000000011;
mem2[548] = 10'b0000000011;
mem2[549] = 10'b0000000011;
mem2[550] = 10'b0000000011;
mem2[551] = 10'b0000000011;
mem2[552] = 10'b0000000011;
mem2[553] = 10'b0000000011;
mem2[554] = 10'b0000000011;
mem2[555] = 10'b0000000011;
mem2[556] = 10'b0000000011;
mem2[557] = 10'b0000000011;
mem2[558] = 10'b0000000011;
mem2[559] = 10'b0000000011;
mem2[560] = 10'b0000000011;
mem2[561] = 10'b0000000011;
mem2[562] = 10'b0000000011;
mem2[563] = 10'b0000000011;
mem2[564] = 10'b0000000011;
mem2[565] = 10'b0000000011;
mem2[566] = 10'b0000000011;
mem2[567] = 10'b0000000011;
mem2[568] = 10'b0000000011;
mem2[569] = 10'b0000000011;
mem2[570] = 10'b0000000011;
mem2[571] = 10'b0000000011;
mem2[572] = 10'b0000000011;
mem2[573] = 10'b0000000011;
mem2[574] = 10'b0000000011;
mem2[575] = 10'b0000000011;
mem2[576] = 10'b0000000011;
mem2[577] = 10'b0000000011;
mem2[578] = 10'b0000000011;
mem2[579] = 10'b0000000011;
mem2[580] = 10'b0000000011;
mem2[581] = 10'b0000000011;
mem2[582] = 10'b0000000011;
mem2[583] = 10'b0000000011;
mem2[584] = 10'b0000000011;
mem2[585] = 10'b0000000011;
mem2[586] = 10'b0000000011;
mem2[587] = 10'b0000000011;
mem2[588] = 10'b0000000011;
mem2[589] = 10'b0000000011;
mem2[590] = 10'b0000000011;
mem2[591] = 10'b0000000011;
mem2[592] = 10'b0000000011;
mem2[593] = 10'b0000000011;
mem2[594] = 10'b0000000011;
mem2[595] = 10'b0000000011;
mem2[596] = 10'b0000000011;
mem2[597] = 10'b0000000011;
mem2[598] = 10'b0000000011;
mem2[599] = 10'b0000000011;
mem2[600] = 10'b0000000011;
mem2[601] = 10'b0000000011;
mem2[602] = 10'b0000000011;
mem2[603] = 10'b0000000011;
mem2[604] = 10'b0000000011;
mem2[605] = 10'b0000000011;
mem2[606] = 10'b0000000011;
mem2[607] = 10'b0000000011;
mem2[608] = 10'b0000000011;
mem2[609] = 10'b0000000011;
mem2[610] = 10'b0000000011;
mem2[611] = 10'b0000000011;
mem2[612] = 10'b0000000100;
mem2[613] = 10'b0000000100;
mem2[614] = 10'b0000000100;
mem2[615] = 10'b0000000100;
mem2[616] = 10'b0000000100;
mem2[617] = 10'b0000000100;
mem2[618] = 10'b0000000100;
mem2[619] = 10'b0000000100;
mem2[620] = 10'b0000000100;
mem2[621] = 10'b0000000100;
mem2[622] = 10'b0000000100;
mem2[623] = 10'b0000000100;
mem2[624] = 10'b0000000100;
mem2[625] = 10'b0000000100;
mem2[626] = 10'b0000000100;
mem2[627] = 10'b0000000100;
mem2[628] = 10'b0000000100;
mem2[629] = 10'b0000000100;
mem2[630] = 10'b0000000100;
mem2[631] = 10'b0000000100;
mem2[632] = 10'b0000000100;
mem2[633] = 10'b0000000100;
mem2[634] = 10'b0000000100;
mem2[635] = 10'b0000000100;
mem2[636] = 10'b0000000100;
mem2[637] = 10'b0000000100;
mem2[638] = 10'b0000000100;
mem2[639] = 10'b0000000100;
mem2[640] = 10'b0000000100;
mem2[641] = 10'b0000000100;
mem2[642] = 10'b0000000100;
mem2[643] = 10'b0000000100;
mem2[644] = 10'b0000000100;
mem2[645] = 10'b0000000100;
mem2[646] = 10'b0000000100;
mem2[647] = 10'b0000000100;
mem2[648] = 10'b0000000100;
mem2[649] = 10'b0000000100;
mem2[650] = 10'b0000000100;
mem2[651] = 10'b0000000100;
mem2[652] = 10'b0000000100;
mem2[653] = 10'b0000000100;
mem2[654] = 10'b0000000100;
mem2[655] = 10'b0000000100;
mem2[656] = 10'b0000000100;
mem2[657] = 10'b0000000100;
mem2[658] = 10'b0000000100;
mem2[659] = 10'b0000000100;
mem2[660] = 10'b0000000100;
mem2[661] = 10'b0000000100;
mem2[662] = 10'b0000000100;
mem2[663] = 10'b0000000100;
mem2[664] = 10'b0000000100;
mem2[665] = 10'b0000000100;
mem2[666] = 10'b0000000100;
mem2[667] = 10'b0000000100;
mem2[668] = 10'b0000000100;
mem2[669] = 10'b0000000100;
mem2[670] = 10'b0000000100;
mem2[671] = 10'b0000000100;
mem2[672] = 10'b0000000100;
mem2[673] = 10'b0000000100;
mem2[674] = 10'b0000000100;
mem2[675] = 10'b0000000100;
mem2[676] = 10'b0000000100;
mem2[677] = 10'b0000000100;
mem2[678] = 10'b0000000100;
mem2[679] = 10'b0000000100;
mem2[680] = 10'b0000000100;
mem2[681] = 10'b0000000100;
mem2[682] = 10'b0000000100;
mem2[683] = 10'b0000000100;
mem2[684] = 10'b0000000101;
mem2[685] = 10'b0000000101;
mem2[686] = 10'b0000000101;
mem2[687] = 10'b0000000101;
mem2[688] = 10'b0000000101;
mem2[689] = 10'b0000000101;
mem2[690] = 10'b0000000101;
mem2[691] = 10'b0000000101;
mem2[692] = 10'b0000000101;
mem2[693] = 10'b0000000101;
mem2[694] = 10'b0000000101;
mem2[695] = 10'b0000000101;
mem2[696] = 10'b0000000101;
mem2[697] = 10'b0000000101;
mem2[698] = 10'b0000000101;
mem2[699] = 10'b0000000101;
mem2[700] = 10'b0000000101;
mem2[701] = 10'b0000000101;
mem2[702] = 10'b0000000101;
mem2[703] = 10'b0000000101;
mem2[704] = 10'b0000000101;
mem2[705] = 10'b0000000101;
mem2[706] = 10'b0000000101;
mem2[707] = 10'b0000000101;
mem2[708] = 10'b0000000101;
mem2[709] = 10'b0000000101;
mem2[710] = 10'b0000000101;
mem2[711] = 10'b0000000101;
mem2[712] = 10'b0000000101;
mem2[713] = 10'b0000000101;
mem2[714] = 10'b0000000101;
mem2[715] = 10'b0000000101;
mem2[716] = 10'b0000000101;
mem2[717] = 10'b0000000101;
mem2[718] = 10'b0000000101;
mem2[719] = 10'b0000000101;
mem2[720] = 10'b0000000101;
mem2[721] = 10'b0000000101;
mem2[722] = 10'b0000000101;
mem2[723] = 10'b0000000101;
mem2[724] = 10'b0000000101;
mem2[725] = 10'b0000000101;
mem2[726] = 10'b0000000101;
mem2[727] = 10'b0000000101;
mem2[728] = 10'b0000000101;
mem2[729] = 10'b0000000101;
mem2[730] = 10'b0000000101;
mem2[731] = 10'b0000000101;
mem2[732] = 10'b0000000101;
mem2[733] = 10'b0000000101;
mem2[734] = 10'b0000000101;
mem2[735] = 10'b0000000101;
mem2[736] = 10'b0000000101;
mem2[737] = 10'b0000000101;
mem2[738] = 10'b0000000101;
mem2[739] = 10'b0000000101;
mem2[740] = 10'b0000000101;
mem2[741] = 10'b0000000101;
mem2[742] = 10'b0000000101;
mem2[743] = 10'b0000000101;
mem2[744] = 10'b0000000101;
mem2[745] = 10'b0000000101;
mem2[746] = 10'b0000000101;
mem2[747] = 10'b0000000101;
mem2[748] = 10'b0000000101;
mem2[749] = 10'b0000000110;
mem2[750] = 10'b0000000110;
mem2[751] = 10'b0000000110;
mem2[752] = 10'b0000000110;
mem2[753] = 10'b0000000110;
mem2[754] = 10'b0000000110;
mem2[755] = 10'b0000000110;
mem2[756] = 10'b0000000110;
mem2[757] = 10'b0000000110;
mem2[758] = 10'b0000000110;
mem2[759] = 10'b0000000110;
mem2[760] = 10'b0000000110;
mem2[761] = 10'b0000000110;
mem2[762] = 10'b0000000110;
mem2[763] = 10'b0000000110;
mem2[764] = 10'b0000000110;
mem2[765] = 10'b0000000110;
mem2[766] = 10'b0000000110;
mem2[767] = 10'b0000000110;
mem2[768] = 10'b0000000110;
mem2[769] = 10'b0000000110;
mem2[770] = 10'b0000000110;
mem2[771] = 10'b0000000110;
mem2[772] = 10'b0000000110;
mem2[773] = 10'b0000000110;
mem2[774] = 10'b0000000110;
mem2[775] = 10'b0000000110;
mem2[776] = 10'b0000000110;
mem2[777] = 10'b0000000110;
mem2[778] = 10'b0000000110;
mem2[779] = 10'b0000000110;
mem2[780] = 10'b0000000110;
mem2[781] = 10'b0000000110;
mem2[782] = 10'b0000000110;
mem2[783] = 10'b0000000110;
mem2[784] = 10'b0000000110;
mem2[785] = 10'b0000000110;
mem2[786] = 10'b0000000110;
mem2[787] = 10'b0000000110;
mem2[788] = 10'b0000000110;
mem2[789] = 10'b0000000110;
mem2[790] = 10'b0000000110;
mem2[791] = 10'b0000000110;
mem2[792] = 10'b0000000110;
mem2[793] = 10'b0000000110;
mem2[794] = 10'b0000000110;
mem2[795] = 10'b0000000110;
mem2[796] = 10'b0000000110;
mem2[797] = 10'b0000000110;
mem2[798] = 10'b0000000110;
mem2[799] = 10'b0000000110;
mem2[800] = 10'b0000000110;
mem2[801] = 10'b0000000110;
mem2[802] = 10'b0000000110;
mem2[803] = 10'b0000000110;
mem2[804] = 10'b0000000110;
mem2[805] = 10'b0000000110;
mem2[806] = 10'b0000000110;
mem2[807] = 10'b0000000110;
mem2[808] = 10'b0000000110;
mem2[809] = 10'b0000000110;
mem2[810] = 10'b0000000111;
mem2[811] = 10'b0000000111;
mem2[812] = 10'b0000000111;
mem2[813] = 10'b0000000111;
mem2[814] = 10'b0000000111;
mem2[815] = 10'b0000000111;
mem2[816] = 10'b0000000111;
mem2[817] = 10'b0000000111;
mem2[818] = 10'b0000000111;
mem2[819] = 10'b0000000111;
mem2[820] = 10'b0000000111;
mem2[821] = 10'b0000000111;
mem2[822] = 10'b0000000111;
mem2[823] = 10'b0000000111;
mem2[824] = 10'b0000000111;
mem2[825] = 10'b0000000111;
mem2[826] = 10'b0000000111;
mem2[827] = 10'b0000000111;
mem2[828] = 10'b0000000111;
mem2[829] = 10'b0000000111;
mem2[830] = 10'b0000000111;
mem2[831] = 10'b0000000111;
mem2[832] = 10'b0000000111;
mem2[833] = 10'b0000000111;
mem2[834] = 10'b0000000111;
mem2[835] = 10'b0000000111;
mem2[836] = 10'b0000000111;
mem2[837] = 10'b0000000111;
mem2[838] = 10'b0000000111;
mem2[839] = 10'b0000000111;
mem2[840] = 10'b0000000111;
mem2[841] = 10'b0000000111;
mem2[842] = 10'b0000000111;
mem2[843] = 10'b0000000111;
mem2[844] = 10'b0000000111;
mem2[845] = 10'b0000000111;
mem2[846] = 10'b0000000111;
mem2[847] = 10'b0000000111;
mem2[848] = 10'b0000000111;
mem2[849] = 10'b0000000111;
mem2[850] = 10'b0000000111;
mem2[851] = 10'b0000000111;
mem2[852] = 10'b0000000111;
mem2[853] = 10'b0000000111;
mem2[854] = 10'b0000000111;
mem2[855] = 10'b0000000111;
mem2[856] = 10'b0000000111;
mem2[857] = 10'b0000000111;
mem2[858] = 10'b0000000111;
mem2[859] = 10'b0000000111;
mem2[860] = 10'b0000000111;
mem2[861] = 10'b0000000111;
mem2[862] = 10'b0000000111;
mem2[863] = 10'b0000000111;
mem2[864] = 10'b0000000111;
mem2[865] = 10'b0000000111;
mem2[866] = 10'b0000001000;
mem2[867] = 10'b0000001000;
mem2[868] = 10'b0000001000;
mem2[869] = 10'b0000001000;
mem2[870] = 10'b0000001000;
mem2[871] = 10'b0000001000;
mem2[872] = 10'b0000001000;
mem2[873] = 10'b0000001000;
mem2[874] = 10'b0000001000;
mem2[875] = 10'b0000001000;
mem2[876] = 10'b0000001000;
mem2[877] = 10'b0000001000;
mem2[878] = 10'b0000001000;
mem2[879] = 10'b0000001000;
mem2[880] = 10'b0000001000;
mem2[881] = 10'b0000001000;
mem2[882] = 10'b0000001000;
mem2[883] = 10'b0000001000;
mem2[884] = 10'b0000001000;
mem2[885] = 10'b0000001000;
mem2[886] = 10'b0000001000;
mem2[887] = 10'b0000001000;
mem2[888] = 10'b0000001000;
mem2[889] = 10'b0000001000;
mem2[890] = 10'b0000001000;
mem2[891] = 10'b0000001000;
mem2[892] = 10'b0000001000;
mem2[893] = 10'b0000001000;
mem2[894] = 10'b0000001000;
mem2[895] = 10'b0000001000;
mem2[896] = 10'b0000001000;
mem2[897] = 10'b0000001000;
mem2[898] = 10'b0000001000;
mem2[899] = 10'b0000001000;
mem2[900] = 10'b0000001000;
mem2[901] = 10'b0000001000;
mem2[902] = 10'b0000001000;
mem2[903] = 10'b0000001000;
mem2[904] = 10'b0000001000;
mem2[905] = 10'b0000001000;
mem2[906] = 10'b0000001000;
mem2[907] = 10'b0000001000;
mem2[908] = 10'b0000001000;
mem2[909] = 10'b0000001000;
mem2[910] = 10'b0000001000;
mem2[911] = 10'b0000001000;
mem2[912] = 10'b0000001000;
mem2[913] = 10'b0000001000;
mem2[914] = 10'b0000001000;
mem2[915] = 10'b0000001000;
mem2[916] = 10'b0000001000;
mem2[917] = 10'b0000001000;
mem2[918] = 10'b0000001001;
mem2[919] = 10'b0000001001;
mem2[920] = 10'b0000001001;
mem2[921] = 10'b0000001001;
mem2[922] = 10'b0000001001;
mem2[923] = 10'b0000001001;
mem2[924] = 10'b0000001001;
mem2[925] = 10'b0000001001;
mem2[926] = 10'b0000001001;
mem2[927] = 10'b0000001001;
mem2[928] = 10'b0000001001;
mem2[929] = 10'b0000001001;
mem2[930] = 10'b0000001001;
mem2[931] = 10'b0000001001;
mem2[932] = 10'b0000001001;
mem2[933] = 10'b0000001001;
mem2[934] = 10'b0000001001;
mem2[935] = 10'b0000001001;
mem2[936] = 10'b0000001001;
mem2[937] = 10'b0000001001;
mem2[938] = 10'b0000001001;
mem2[939] = 10'b0000001001;
mem2[940] = 10'b0000001001;
mem2[941] = 10'b0000001001;
mem2[942] = 10'b0000001001;
mem2[943] = 10'b0000001001;
mem2[944] = 10'b0000001001;
mem2[945] = 10'b0000001001;
mem2[946] = 10'b0000001001;
mem2[947] = 10'b0000001001;
mem2[948] = 10'b0000001001;
mem2[949] = 10'b0000001001;
mem2[950] = 10'b0000001001;
mem2[951] = 10'b0000001001;
mem2[952] = 10'b0000001001;
mem2[953] = 10'b0000001001;
mem2[954] = 10'b0000001001;
mem2[955] = 10'b0000001001;
mem2[956] = 10'b0000001001;
mem2[957] = 10'b0000001001;
mem2[958] = 10'b0000001001;
mem2[959] = 10'b0000001001;
mem2[960] = 10'b0000001001;
mem2[961] = 10'b0000001001;
mem2[962] = 10'b0000001001;
mem2[963] = 10'b0000001001;
mem2[964] = 10'b0000001001;
mem2[965] = 10'b0000001001;
mem2[966] = 10'b0000001001;
mem2[967] = 10'b0000001001;
mem2[968] = 10'b0000001010;
mem2[969] = 10'b0000001010;
mem2[970] = 10'b0000001010;
mem2[971] = 10'b0000001010;
mem2[972] = 10'b0000001010;
mem2[973] = 10'b0000001010;
mem2[974] = 10'b0000001010;
mem2[975] = 10'b0000001010;
mem2[976] = 10'b0000001010;
mem2[977] = 10'b0000001010;
mem2[978] = 10'b0000001010;
mem2[979] = 10'b0000001010;
mem2[980] = 10'b0000001010;
mem2[981] = 10'b0000001010;
mem2[982] = 10'b0000001010;
mem2[983] = 10'b0000001010;
mem2[984] = 10'b0000001010;
mem2[985] = 10'b0000001010;
mem2[986] = 10'b0000001010;
mem2[987] = 10'b0000001010;
mem2[988] = 10'b0000001010;
mem2[989] = 10'b0000001010;
mem2[990] = 10'b0000001010;
mem2[991] = 10'b0000001010;
mem2[992] = 10'b0000001010;
mem2[993] = 10'b0000001010;
mem2[994] = 10'b0000001010;
mem2[995] = 10'b0000001010;
mem2[996] = 10'b0000001010;
mem2[997] = 10'b0000001010;
mem2[998] = 10'b0000001010;
mem2[999] = 10'b0000001010;
mem2[1000] = 10'b0000001010;
mem2[1001] = 10'b0000001010;
mem2[1002] = 10'b0000001010;
mem2[1003] = 10'b0000001010;
mem2[1004] = 10'b0000001010;
mem2[1005] = 10'b0000001010;
mem2[1006] = 10'b0000001010;
mem2[1007] = 10'b0000001010;
mem2[1008] = 10'b0000001010;
mem2[1009] = 10'b0000001010;
mem2[1010] = 10'b0000001010;
mem2[1011] = 10'b0000001010;
mem2[1012] = 10'b0000001010;
mem2[1013] = 10'b0000001010;
mem2[1014] = 10'b0000001010;
mem2[1015] = 10'b0000001010;
mem2[1016] = 10'b0000001011;
mem2[1017] = 10'b0000001011;
mem2[1018] = 10'b0000001011;
mem2[1019] = 10'b0000001011;
mem2[1020] = 10'b0000001011;
mem2[1021] = 10'b0000001011;
mem2[1022] = 10'b0000001011;
mem2[1023] = 10'b0000001011;
mem2[1024] = 10'b0000001011;
mem2[1025] = 10'b0000001011;
mem2[1026] = 10'b0000001011;
mem2[1027] = 10'b0000001011;
mem2[1028] = 10'b0000001011;
mem2[1029] = 10'b0000001011;
mem2[1030] = 10'b0000001011;
mem2[1031] = 10'b0000001011;
mem2[1032] = 10'b0000001011;
mem2[1033] = 10'b0000001011;
mem2[1034] = 10'b0000001011;
mem2[1035] = 10'b0000001011;
mem2[1036] = 10'b0000001011;
mem2[1037] = 10'b0000001011;
mem2[1038] = 10'b0000001011;
mem2[1039] = 10'b0000001011;
mem2[1040] = 10'b0000001011;
mem2[1041] = 10'b0000001011;
mem2[1042] = 10'b0000001011;
mem2[1043] = 10'b0000001011;
mem2[1044] = 10'b0000001011;
mem2[1045] = 10'b0000001011;
mem2[1046] = 10'b0000001011;
mem2[1047] = 10'b0000001011;
mem2[1048] = 10'b0000001011;
mem2[1049] = 10'b0000001011;
mem2[1050] = 10'b0000001011;
mem2[1051] = 10'b0000001011;
mem2[1052] = 10'b0000001011;
mem2[1053] = 10'b0000001011;
mem2[1054] = 10'b0000001011;
mem2[1055] = 10'b0000001011;
mem2[1056] = 10'b0000001011;
mem2[1057] = 10'b0000001011;
mem2[1058] = 10'b0000001011;
mem2[1059] = 10'b0000001011;
mem2[1060] = 10'b0000001011;
mem2[1061] = 10'b0000001100;
mem2[1062] = 10'b0000001100;
mem2[1063] = 10'b0000001100;
mem2[1064] = 10'b0000001100;
mem2[1065] = 10'b0000001100;
mem2[1066] = 10'b0000001100;
mem2[1067] = 10'b0000001100;
mem2[1068] = 10'b0000001100;
mem2[1069] = 10'b0000001100;
mem2[1070] = 10'b0000001100;
mem2[1071] = 10'b0000001100;
mem2[1072] = 10'b0000001100;
mem2[1073] = 10'b0000001100;
mem2[1074] = 10'b0000001100;
mem2[1075] = 10'b0000001100;
mem2[1076] = 10'b0000001100;
mem2[1077] = 10'b0000001100;
mem2[1078] = 10'b0000001100;
mem2[1079] = 10'b0000001100;
mem2[1080] = 10'b0000001100;
mem2[1081] = 10'b0000001100;
mem2[1082] = 10'b0000001100;
mem2[1083] = 10'b0000001100;
mem2[1084] = 10'b0000001100;
mem2[1085] = 10'b0000001100;
mem2[1086] = 10'b0000001100;
mem2[1087] = 10'b0000001100;
mem2[1088] = 10'b0000001100;
mem2[1089] = 10'b0000001100;
mem2[1090] = 10'b0000001100;
mem2[1091] = 10'b0000001100;
mem2[1092] = 10'b0000001100;
mem2[1093] = 10'b0000001100;
mem2[1094] = 10'b0000001100;
mem2[1095] = 10'b0000001100;
mem2[1096] = 10'b0000001100;
mem2[1097] = 10'b0000001100;
mem2[1098] = 10'b0000001100;
mem2[1099] = 10'b0000001100;
mem2[1100] = 10'b0000001100;
mem2[1101] = 10'b0000001100;
mem2[1102] = 10'b0000001100;
mem2[1103] = 10'b0000001100;
mem2[1104] = 10'b0000001101;
mem2[1105] = 10'b0000001101;
mem2[1106] = 10'b0000001101;
mem2[1107] = 10'b0000001101;
mem2[1108] = 10'b0000001101;
mem2[1109] = 10'b0000001101;
mem2[1110] = 10'b0000001101;
mem2[1111] = 10'b0000001101;
mem2[1112] = 10'b0000001101;
mem2[1113] = 10'b0000001101;
mem2[1114] = 10'b0000001101;
mem2[1115] = 10'b0000001101;
mem2[1116] = 10'b0000001101;
mem2[1117] = 10'b0000001101;
mem2[1118] = 10'b0000001101;
mem2[1119] = 10'b0000001101;
mem2[1120] = 10'b0000001101;
mem2[1121] = 10'b0000001101;
mem2[1122] = 10'b0000001101;
mem2[1123] = 10'b0000001101;
mem2[1124] = 10'b0000001101;
mem2[1125] = 10'b0000001101;
mem2[1126] = 10'b0000001101;
mem2[1127] = 10'b0000001101;
mem2[1128] = 10'b0000001101;
mem2[1129] = 10'b0000001101;
mem2[1130] = 10'b0000001101;
mem2[1131] = 10'b0000001101;
mem2[1132] = 10'b0000001101;
mem2[1133] = 10'b0000001101;
mem2[1134] = 10'b0000001101;
mem2[1135] = 10'b0000001101;
mem2[1136] = 10'b0000001101;
mem2[1137] = 10'b0000001101;
mem2[1138] = 10'b0000001101;
mem2[1139] = 10'b0000001101;
mem2[1140] = 10'b0000001101;
mem2[1141] = 10'b0000001101;
mem2[1142] = 10'b0000001101;
mem2[1143] = 10'b0000001101;
mem2[1144] = 10'b0000001101;
mem2[1145] = 10'b0000001101;
mem2[1146] = 10'b0000001110;
mem2[1147] = 10'b0000001110;
mem2[1148] = 10'b0000001110;
mem2[1149] = 10'b0000001110;
mem2[1150] = 10'b0000001110;
mem2[1151] = 10'b0000001110;
mem2[1152] = 10'b0000001110;
mem2[1153] = 10'b0000001110;
mem2[1154] = 10'b0000001110;
mem2[1155] = 10'b0000001110;
mem2[1156] = 10'b0000001110;
mem2[1157] = 10'b0000001110;
mem2[1158] = 10'b0000001110;
mem2[1159] = 10'b0000001110;
mem2[1160] = 10'b0000001110;
mem2[1161] = 10'b0000001110;
mem2[1162] = 10'b0000001110;
mem2[1163] = 10'b0000001110;
mem2[1164] = 10'b0000001110;
mem2[1165] = 10'b0000001110;
mem2[1166] = 10'b0000001110;
mem2[1167] = 10'b0000001110;
mem2[1168] = 10'b0000001110;
mem2[1169] = 10'b0000001110;
mem2[1170] = 10'b0000001110;
mem2[1171] = 10'b0000001110;
mem2[1172] = 10'b0000001110;
mem2[1173] = 10'b0000001110;
mem2[1174] = 10'b0000001110;
mem2[1175] = 10'b0000001110;
mem2[1176] = 10'b0000001110;
mem2[1177] = 10'b0000001110;
mem2[1178] = 10'b0000001110;
mem2[1179] = 10'b0000001110;
mem2[1180] = 10'b0000001110;
mem2[1181] = 10'b0000001110;
mem2[1182] = 10'b0000001110;
mem2[1183] = 10'b0000001110;
mem2[1184] = 10'b0000001110;
mem2[1185] = 10'b0000001110;
mem2[1186] = 10'b0000001110;
mem2[1187] = 10'b0000001111;
mem2[1188] = 10'b0000001111;
mem2[1189] = 10'b0000001111;
mem2[1190] = 10'b0000001111;
mem2[1191] = 10'b0000001111;
mem2[1192] = 10'b0000001111;
mem2[1193] = 10'b0000001111;
mem2[1194] = 10'b0000001111;
mem2[1195] = 10'b0000001111;
mem2[1196] = 10'b0000001111;
mem2[1197] = 10'b0000001111;
mem2[1198] = 10'b0000001111;
mem2[1199] = 10'b0000001111;
mem2[1200] = 10'b0000001111;
mem2[1201] = 10'b0000001111;
mem2[1202] = 10'b0000001111;
mem2[1203] = 10'b0000001111;
mem2[1204] = 10'b0000001111;
mem2[1205] = 10'b0000001111;
mem2[1206] = 10'b0000001111;
mem2[1207] = 10'b0000001111;
mem2[1208] = 10'b0000001111;
mem2[1209] = 10'b0000001111;
mem2[1210] = 10'b0000001111;
mem2[1211] = 10'b0000001111;
mem2[1212] = 10'b0000001111;
mem2[1213] = 10'b0000001111;
mem2[1214] = 10'b0000001111;
mem2[1215] = 10'b0000001111;
mem2[1216] = 10'b0000001111;
mem2[1217] = 10'b0000001111;
mem2[1218] = 10'b0000001111;
mem2[1219] = 10'b0000001111;
mem2[1220] = 10'b0000001111;
mem2[1221] = 10'b0000001111;
mem2[1222] = 10'b0000001111;
mem2[1223] = 10'b0000001111;
mem2[1224] = 10'b0000001111;
mem2[1225] = 10'b0000001111;
mem2[1226] = 10'b0000010000;
mem2[1227] = 10'b0000010000;
mem2[1228] = 10'b0000010000;
mem2[1229] = 10'b0000010000;
mem2[1230] = 10'b0000010000;
mem2[1231] = 10'b0000010000;
mem2[1232] = 10'b0000010000;
mem2[1233] = 10'b0000010000;
mem2[1234] = 10'b0000010000;
mem2[1235] = 10'b0000010000;
mem2[1236] = 10'b0000010000;
mem2[1237] = 10'b0000010000;
mem2[1238] = 10'b0000010000;
mem2[1239] = 10'b0000010000;
mem2[1240] = 10'b0000010000;
mem2[1241] = 10'b0000010000;
mem2[1242] = 10'b0000010000;
mem2[1243] = 10'b0000010000;
mem2[1244] = 10'b0000010000;
mem2[1245] = 10'b0000010000;
mem2[1246] = 10'b0000010000;
mem2[1247] = 10'b0000010000;
mem2[1248] = 10'b0000010000;
mem2[1249] = 10'b0000010000;
mem2[1250] = 10'b0000010000;
mem2[1251] = 10'b0000010000;
mem2[1252] = 10'b0000010000;
mem2[1253] = 10'b0000010000;
mem2[1254] = 10'b0000010000;
mem2[1255] = 10'b0000010000;
mem2[1256] = 10'b0000010000;
mem2[1257] = 10'b0000010000;
mem2[1258] = 10'b0000010000;
mem2[1259] = 10'b0000010000;
mem2[1260] = 10'b0000010000;
mem2[1261] = 10'b0000010000;
mem2[1262] = 10'b0000010000;
mem2[1263] = 10'b0000010000;
mem2[1264] = 10'b0000010001;
mem2[1265] = 10'b0000010001;
mem2[1266] = 10'b0000010001;
mem2[1267] = 10'b0000010001;
mem2[1268] = 10'b0000010001;
mem2[1269] = 10'b0000010001;
mem2[1270] = 10'b0000010001;
mem2[1271] = 10'b0000010001;
mem2[1272] = 10'b0000010001;
mem2[1273] = 10'b0000010001;
mem2[1274] = 10'b0000010001;
mem2[1275] = 10'b0000010001;
mem2[1276] = 10'b0000010001;
mem2[1277] = 10'b0000010001;
mem2[1278] = 10'b0000010001;
mem2[1279] = 10'b0000010001;
mem2[1280] = 10'b0000010001;
mem2[1281] = 10'b0000010001;
mem2[1282] = 10'b0000010001;
mem2[1283] = 10'b0000010001;
mem2[1284] = 10'b0000010001;
mem2[1285] = 10'b0000010001;
mem2[1286] = 10'b0000010001;
mem2[1287] = 10'b0000010001;
mem2[1288] = 10'b0000010001;
mem2[1289] = 10'b0000010001;
mem2[1290] = 10'b0000010001;
mem2[1291] = 10'b0000010001;
mem2[1292] = 10'b0000010001;
mem2[1293] = 10'b0000010001;
mem2[1294] = 10'b0000010001;
mem2[1295] = 10'b0000010001;
mem2[1296] = 10'b0000010001;
mem2[1297] = 10'b0000010001;
mem2[1298] = 10'b0000010001;
mem2[1299] = 10'b0000010001;
mem2[1300] = 10'b0000010010;
mem2[1301] = 10'b0000010010;
mem2[1302] = 10'b0000010010;
mem2[1303] = 10'b0000010010;
mem2[1304] = 10'b0000010010;
mem2[1305] = 10'b0000010010;
mem2[1306] = 10'b0000010010;
mem2[1307] = 10'b0000010010;
mem2[1308] = 10'b0000010010;
mem2[1309] = 10'b0000010010;
mem2[1310] = 10'b0000010010;
mem2[1311] = 10'b0000010010;
mem2[1312] = 10'b0000010010;
mem2[1313] = 10'b0000010010;
mem2[1314] = 10'b0000010010;
mem2[1315] = 10'b0000010010;
mem2[1316] = 10'b0000010010;
mem2[1317] = 10'b0000010010;
mem2[1318] = 10'b0000010010;
mem2[1319] = 10'b0000010010;
mem2[1320] = 10'b0000010010;
mem2[1321] = 10'b0000010010;
mem2[1322] = 10'b0000010010;
mem2[1323] = 10'b0000010010;
mem2[1324] = 10'b0000010010;
mem2[1325] = 10'b0000010010;
mem2[1326] = 10'b0000010010;
mem2[1327] = 10'b0000010010;
mem2[1328] = 10'b0000010010;
mem2[1329] = 10'b0000010010;
mem2[1330] = 10'b0000010010;
mem2[1331] = 10'b0000010010;
mem2[1332] = 10'b0000010010;
mem2[1333] = 10'b0000010010;
mem2[1334] = 10'b0000010010;
mem2[1335] = 10'b0000010010;
mem2[1336] = 10'b0000010011;
mem2[1337] = 10'b0000010011;
mem2[1338] = 10'b0000010011;
mem2[1339] = 10'b0000010011;
mem2[1340] = 10'b0000010011;
mem2[1341] = 10'b0000010011;
mem2[1342] = 10'b0000010011;
mem2[1343] = 10'b0000010011;
mem2[1344] = 10'b0000010011;
mem2[1345] = 10'b0000010011;
mem2[1346] = 10'b0000010011;
mem2[1347] = 10'b0000010011;
mem2[1348] = 10'b0000010011;
mem2[1349] = 10'b0000010011;
mem2[1350] = 10'b0000010011;
mem2[1351] = 10'b0000010011;
mem2[1352] = 10'b0000010011;
mem2[1353] = 10'b0000010011;
mem2[1354] = 10'b0000010011;
mem2[1355] = 10'b0000010011;
mem2[1356] = 10'b0000010011;
mem2[1357] = 10'b0000010011;
mem2[1358] = 10'b0000010011;
mem2[1359] = 10'b0000010011;
mem2[1360] = 10'b0000010011;
mem2[1361] = 10'b0000010011;
mem2[1362] = 10'b0000010011;
mem2[1363] = 10'b0000010011;
mem2[1364] = 10'b0000010011;
mem2[1365] = 10'b0000010011;
mem2[1366] = 10'b0000010011;
mem2[1367] = 10'b0000010011;
mem2[1368] = 10'b0000010011;
mem2[1369] = 10'b0000010011;
mem2[1370] = 10'b0000010011;
mem2[1371] = 10'b0000010100;
mem2[1372] = 10'b0000010100;
mem2[1373] = 10'b0000010100;
mem2[1374] = 10'b0000010100;
mem2[1375] = 10'b0000010100;
mem2[1376] = 10'b0000010100;
mem2[1377] = 10'b0000010100;
mem2[1378] = 10'b0000010100;
mem2[1379] = 10'b0000010100;
mem2[1380] = 10'b0000010100;
mem2[1381] = 10'b0000010100;
mem2[1382] = 10'b0000010100;
mem2[1383] = 10'b0000010100;
mem2[1384] = 10'b0000010100;
mem2[1385] = 10'b0000010100;
mem2[1386] = 10'b0000010100;
mem2[1387] = 10'b0000010100;
mem2[1388] = 10'b0000010100;
mem2[1389] = 10'b0000010100;
mem2[1390] = 10'b0000010100;
mem2[1391] = 10'b0000010100;
mem2[1392] = 10'b0000010100;
mem2[1393] = 10'b0000010100;
mem2[1394] = 10'b0000010100;
mem2[1395] = 10'b0000010100;
mem2[1396] = 10'b0000010100;
mem2[1397] = 10'b0000010100;
mem2[1398] = 10'b0000010100;
mem2[1399] = 10'b0000010100;
mem2[1400] = 10'b0000010100;
mem2[1401] = 10'b0000010100;
mem2[1402] = 10'b0000010100;
mem2[1403] = 10'b0000010100;
mem2[1404] = 10'b0000010100;
mem2[1405] = 10'b0000010101;
mem2[1406] = 10'b0000010101;
mem2[1407] = 10'b0000010101;
mem2[1408] = 10'b0000010101;
mem2[1409] = 10'b0000010101;
mem2[1410] = 10'b0000010101;
mem2[1411] = 10'b0000010101;
mem2[1412] = 10'b0000010101;
mem2[1413] = 10'b0000010101;
mem2[1414] = 10'b0000010101;
mem2[1415] = 10'b0000010101;
mem2[1416] = 10'b0000010101;
mem2[1417] = 10'b0000010101;
mem2[1418] = 10'b0000010101;
mem2[1419] = 10'b0000010101;
mem2[1420] = 10'b0000010101;
mem2[1421] = 10'b0000010101;
mem2[1422] = 10'b0000010101;
mem2[1423] = 10'b0000010101;
mem2[1424] = 10'b0000010101;
mem2[1425] = 10'b0000010101;
mem2[1426] = 10'b0000010101;
mem2[1427] = 10'b0000010101;
mem2[1428] = 10'b0000010101;
mem2[1429] = 10'b0000010101;
mem2[1430] = 10'b0000010101;
mem2[1431] = 10'b0000010101;
mem2[1432] = 10'b0000010101;
mem2[1433] = 10'b0000010101;
mem2[1434] = 10'b0000010101;
mem2[1435] = 10'b0000010101;
mem2[1436] = 10'b0000010101;
mem2[1437] = 10'b0000010101;
mem2[1438] = 10'b0000010101;
mem2[1439] = 10'b0000010110;
mem2[1440] = 10'b0000010110;
mem2[1441] = 10'b0000010110;
mem2[1442] = 10'b0000010110;
mem2[1443] = 10'b0000010110;
mem2[1444] = 10'b0000010110;
mem2[1445] = 10'b0000010110;
mem2[1446] = 10'b0000010110;
mem2[1447] = 10'b0000010110;
mem2[1448] = 10'b0000010110;
mem2[1449] = 10'b0000010110;
mem2[1450] = 10'b0000010110;
mem2[1451] = 10'b0000010110;
mem2[1452] = 10'b0000010110;
mem2[1453] = 10'b0000010110;
mem2[1454] = 10'b0000010110;
mem2[1455] = 10'b0000010110;
mem2[1456] = 10'b0000010110;
mem2[1457] = 10'b0000010110;
mem2[1458] = 10'b0000010110;
mem2[1459] = 10'b0000010110;
mem2[1460] = 10'b0000010110;
mem2[1461] = 10'b0000010110;
mem2[1462] = 10'b0000010110;
mem2[1463] = 10'b0000010110;
mem2[1464] = 10'b0000010110;
mem2[1465] = 10'b0000010110;
mem2[1466] = 10'b0000010110;
mem2[1467] = 10'b0000010110;
mem2[1468] = 10'b0000010110;
mem2[1469] = 10'b0000010110;
mem2[1470] = 10'b0000010110;
mem2[1471] = 10'b0000010111;
mem2[1472] = 10'b0000010111;
mem2[1473] = 10'b0000010111;
mem2[1474] = 10'b0000010111;
mem2[1475] = 10'b0000010111;
mem2[1476] = 10'b0000010111;
mem2[1477] = 10'b0000010111;
mem2[1478] = 10'b0000010111;
mem2[1479] = 10'b0000010111;
mem2[1480] = 10'b0000010111;
mem2[1481] = 10'b0000010111;
mem2[1482] = 10'b0000010111;
mem2[1483] = 10'b0000010111;
mem2[1484] = 10'b0000010111;
mem2[1485] = 10'b0000010111;
mem2[1486] = 10'b0000010111;
mem2[1487] = 10'b0000010111;
mem2[1488] = 10'b0000010111;
mem2[1489] = 10'b0000010111;
mem2[1490] = 10'b0000010111;
mem2[1491] = 10'b0000010111;
mem2[1492] = 10'b0000010111;
mem2[1493] = 10'b0000010111;
mem2[1494] = 10'b0000010111;
mem2[1495] = 10'b0000010111;
mem2[1496] = 10'b0000010111;
mem2[1497] = 10'b0000010111;
mem2[1498] = 10'b0000010111;
mem2[1499] = 10'b0000010111;
mem2[1500] = 10'b0000010111;
mem2[1501] = 10'b0000010111;
mem2[1502] = 10'b0000010111;
mem2[1503] = 10'b0000011000;
mem2[1504] = 10'b0000011000;
mem2[1505] = 10'b0000011000;
mem2[1506] = 10'b0000011000;
mem2[1507] = 10'b0000011000;
mem2[1508] = 10'b0000011000;
mem2[1509] = 10'b0000011000;
mem2[1510] = 10'b0000011000;
mem2[1511] = 10'b0000011000;
mem2[1512] = 10'b0000011000;
mem2[1513] = 10'b0000011000;
mem2[1514] = 10'b0000011000;
mem2[1515] = 10'b0000011000;
mem2[1516] = 10'b0000011000;
mem2[1517] = 10'b0000011000;
mem2[1518] = 10'b0000011000;
mem2[1519] = 10'b0000011000;
mem2[1520] = 10'b0000011000;
mem2[1521] = 10'b0000011000;
mem2[1522] = 10'b0000011000;
mem2[1523] = 10'b0000011000;
mem2[1524] = 10'b0000011000;
mem2[1525] = 10'b0000011000;
mem2[1526] = 10'b0000011000;
mem2[1527] = 10'b0000011000;
mem2[1528] = 10'b0000011000;
mem2[1529] = 10'b0000011000;
mem2[1530] = 10'b0000011000;
mem2[1531] = 10'b0000011000;
mem2[1532] = 10'b0000011000;
mem2[1533] = 10'b0000011000;
mem2[1534] = 10'b0000011001;
mem2[1535] = 10'b0000011001;
mem2[1536] = 10'b0000011001;
mem2[1537] = 10'b0000011001;
mem2[1538] = 10'b0000011001;
mem2[1539] = 10'b0000011001;
mem2[1540] = 10'b0000011001;
mem2[1541] = 10'b0000011001;
mem2[1542] = 10'b0000011001;
mem2[1543] = 10'b0000011001;
mem2[1544] = 10'b0000011001;
mem2[1545] = 10'b0000011001;
mem2[1546] = 10'b0000011001;
mem2[1547] = 10'b0000011001;
mem2[1548] = 10'b0000011001;
mem2[1549] = 10'b0000011001;
mem2[1550] = 10'b0000011001;
mem2[1551] = 10'b0000011001;
mem2[1552] = 10'b0000011001;
mem2[1553] = 10'b0000011001;
mem2[1554] = 10'b0000011001;
mem2[1555] = 10'b0000011001;
mem2[1556] = 10'b0000011001;
mem2[1557] = 10'b0000011001;
mem2[1558] = 10'b0000011001;
mem2[1559] = 10'b0000011001;
mem2[1560] = 10'b0000011001;
mem2[1561] = 10'b0000011001;
mem2[1562] = 10'b0000011001;
mem2[1563] = 10'b0000011001;
mem2[1564] = 10'b0000011001;
mem2[1565] = 10'b0000011010;
mem2[1566] = 10'b0000011010;
mem2[1567] = 10'b0000011010;
mem2[1568] = 10'b0000011010;
mem2[1569] = 10'b0000011010;
mem2[1570] = 10'b0000011010;
mem2[1571] = 10'b0000011010;
mem2[1572] = 10'b0000011010;
mem2[1573] = 10'b0000011010;
mem2[1574] = 10'b0000011010;
mem2[1575] = 10'b0000011010;
mem2[1576] = 10'b0000011010;
mem2[1577] = 10'b0000011010;
mem2[1578] = 10'b0000011010;
mem2[1579] = 10'b0000011010;
mem2[1580] = 10'b0000011010;
mem2[1581] = 10'b0000011010;
mem2[1582] = 10'b0000011010;
mem2[1583] = 10'b0000011010;
mem2[1584] = 10'b0000011010;
mem2[1585] = 10'b0000011010;
mem2[1586] = 10'b0000011010;
mem2[1587] = 10'b0000011010;
mem2[1588] = 10'b0000011010;
mem2[1589] = 10'b0000011010;
mem2[1590] = 10'b0000011010;
mem2[1591] = 10'b0000011010;
mem2[1592] = 10'b0000011010;
mem2[1593] = 10'b0000011010;
mem2[1594] = 10'b0000011010;
mem2[1595] = 10'b0000011011;
mem2[1596] = 10'b0000011011;
mem2[1597] = 10'b0000011011;
mem2[1598] = 10'b0000011011;
mem2[1599] = 10'b0000011011;
mem2[1600] = 10'b0000011011;
mem2[1601] = 10'b0000011011;
mem2[1602] = 10'b0000011011;
mem2[1603] = 10'b0000011011;
mem2[1604] = 10'b0000011011;
mem2[1605] = 10'b0000011011;
mem2[1606] = 10'b0000011011;
mem2[1607] = 10'b0000011011;
mem2[1608] = 10'b0000011011;
mem2[1609] = 10'b0000011011;
mem2[1610] = 10'b0000011011;
mem2[1611] = 10'b0000011011;
mem2[1612] = 10'b0000011011;
mem2[1613] = 10'b0000011011;
mem2[1614] = 10'b0000011011;
mem2[1615] = 10'b0000011011;
mem2[1616] = 10'b0000011011;
mem2[1617] = 10'b0000011011;
mem2[1618] = 10'b0000011011;
mem2[1619] = 10'b0000011011;
mem2[1620] = 10'b0000011011;
mem2[1621] = 10'b0000011011;
mem2[1622] = 10'b0000011011;
mem2[1623] = 10'b0000011011;
mem2[1624] = 10'b0000011011;
mem2[1625] = 10'b0000011100;
mem2[1626] = 10'b0000011100;
mem2[1627] = 10'b0000011100;
mem2[1628] = 10'b0000011100;
mem2[1629] = 10'b0000011100;
mem2[1630] = 10'b0000011100;
mem2[1631] = 10'b0000011100;
mem2[1632] = 10'b0000011100;
mem2[1633] = 10'b0000011100;
mem2[1634] = 10'b0000011100;
mem2[1635] = 10'b0000011100;
mem2[1636] = 10'b0000011100;
mem2[1637] = 10'b0000011100;
mem2[1638] = 10'b0000011100;
mem2[1639] = 10'b0000011100;
mem2[1640] = 10'b0000011100;
mem2[1641] = 10'b0000011100;
mem2[1642] = 10'b0000011100;
mem2[1643] = 10'b0000011100;
mem2[1644] = 10'b0000011100;
mem2[1645] = 10'b0000011100;
mem2[1646] = 10'b0000011100;
mem2[1647] = 10'b0000011100;
mem2[1648] = 10'b0000011100;
mem2[1649] = 10'b0000011100;
mem2[1650] = 10'b0000011100;
mem2[1651] = 10'b0000011100;
mem2[1652] = 10'b0000011100;
mem2[1653] = 10'b0000011100;
mem2[1654] = 10'b0000011101;
mem2[1655] = 10'b0000011101;
mem2[1656] = 10'b0000011101;
mem2[1657] = 10'b0000011101;
mem2[1658] = 10'b0000011101;
mem2[1659] = 10'b0000011101;
mem2[1660] = 10'b0000011101;
mem2[1661] = 10'b0000011101;
mem2[1662] = 10'b0000011101;
mem2[1663] = 10'b0000011101;
mem2[1664] = 10'b0000011101;
mem2[1665] = 10'b0000011101;
mem2[1666] = 10'b0000011101;
mem2[1667] = 10'b0000011101;
mem2[1668] = 10'b0000011101;
mem2[1669] = 10'b0000011101;
mem2[1670] = 10'b0000011101;
mem2[1671] = 10'b0000011101;
mem2[1672] = 10'b0000011101;
mem2[1673] = 10'b0000011101;
mem2[1674] = 10'b0000011101;
mem2[1675] = 10'b0000011101;
mem2[1676] = 10'b0000011101;
mem2[1677] = 10'b0000011101;
mem2[1678] = 10'b0000011101;
mem2[1679] = 10'b0000011101;
mem2[1680] = 10'b0000011101;
mem2[1681] = 10'b0000011101;
mem2[1682] = 10'b0000011110;
mem2[1683] = 10'b0000011110;
mem2[1684] = 10'b0000011110;
mem2[1685] = 10'b0000011110;
mem2[1686] = 10'b0000011110;
mem2[1687] = 10'b0000011110;
mem2[1688] = 10'b0000011110;
mem2[1689] = 10'b0000011110;
mem2[1690] = 10'b0000011110;
mem2[1691] = 10'b0000011110;
mem2[1692] = 10'b0000011110;
mem2[1693] = 10'b0000011110;
mem2[1694] = 10'b0000011110;
mem2[1695] = 10'b0000011110;
mem2[1696] = 10'b0000011110;
mem2[1697] = 10'b0000011110;
mem2[1698] = 10'b0000011110;
mem2[1699] = 10'b0000011110;
mem2[1700] = 10'b0000011110;
mem2[1701] = 10'b0000011110;
mem2[1702] = 10'b0000011110;
mem2[1703] = 10'b0000011110;
mem2[1704] = 10'b0000011110;
mem2[1705] = 10'b0000011110;
mem2[1706] = 10'b0000011110;
mem2[1707] = 10'b0000011110;
mem2[1708] = 10'b0000011110;
mem2[1709] = 10'b0000011110;
mem2[1710] = 10'b0000011111;
mem2[1711] = 10'b0000011111;
mem2[1712] = 10'b0000011111;
mem2[1713] = 10'b0000011111;
mem2[1714] = 10'b0000011111;
mem2[1715] = 10'b0000011111;
mem2[1716] = 10'b0000011111;
mem2[1717] = 10'b0000011111;
mem2[1718] = 10'b0000011111;
mem2[1719] = 10'b0000011111;
mem2[1720] = 10'b0000011111;
mem2[1721] = 10'b0000011111;
mem2[1722] = 10'b0000011111;
mem2[1723] = 10'b0000011111;
mem2[1724] = 10'b0000011111;
mem2[1725] = 10'b0000011111;
mem2[1726] = 10'b0000011111;
mem2[1727] = 10'b0000011111;
mem2[1728] = 10'b0000011111;
mem2[1729] = 10'b0000011111;
mem2[1730] = 10'b0000011111;
mem2[1731] = 10'b0000011111;
mem2[1732] = 10'b0000011111;
mem2[1733] = 10'b0000011111;
mem2[1734] = 10'b0000011111;
mem2[1735] = 10'b0000011111;
mem2[1736] = 10'b0000011111;
mem2[1737] = 10'b0000011111;
mem2[1738] = 10'b0000100000;
mem2[1739] = 10'b0000100000;
mem2[1740] = 10'b0000100000;
mem2[1741] = 10'b0000100000;
mem2[1742] = 10'b0000100000;
mem2[1743] = 10'b0000100000;
mem2[1744] = 10'b0000100000;
mem2[1745] = 10'b0000100000;
mem2[1746] = 10'b0000100000;
mem2[1747] = 10'b0000100000;
mem2[1748] = 10'b0000100000;
mem2[1749] = 10'b0000100000;
mem2[1750] = 10'b0000100000;
mem2[1751] = 10'b0000100000;
mem2[1752] = 10'b0000100000;
mem2[1753] = 10'b0000100000;
mem2[1754] = 10'b0000100000;
mem2[1755] = 10'b0000100000;
mem2[1756] = 10'b0000100000;
mem2[1757] = 10'b0000100000;
mem2[1758] = 10'b0000100000;
mem2[1759] = 10'b0000100000;
mem2[1760] = 10'b0000100000;
mem2[1761] = 10'b0000100000;
mem2[1762] = 10'b0000100000;
mem2[1763] = 10'b0000100000;
mem2[1764] = 10'b0000100000;
mem2[1765] = 10'b0000100001;
mem2[1766] = 10'b0000100001;
mem2[1767] = 10'b0000100001;
mem2[1768] = 10'b0000100001;
mem2[1769] = 10'b0000100001;
mem2[1770] = 10'b0000100001;
mem2[1771] = 10'b0000100001;
mem2[1772] = 10'b0000100001;
mem2[1773] = 10'b0000100001;
mem2[1774] = 10'b0000100001;
mem2[1775] = 10'b0000100001;
mem2[1776] = 10'b0000100001;
mem2[1777] = 10'b0000100001;
mem2[1778] = 10'b0000100001;
mem2[1779] = 10'b0000100001;
mem2[1780] = 10'b0000100001;
mem2[1781] = 10'b0000100001;
mem2[1782] = 10'b0000100001;
mem2[1783] = 10'b0000100001;
mem2[1784] = 10'b0000100001;
mem2[1785] = 10'b0000100001;
mem2[1786] = 10'b0000100001;
mem2[1787] = 10'b0000100001;
mem2[1788] = 10'b0000100001;
mem2[1789] = 10'b0000100001;
mem2[1790] = 10'b0000100001;
mem2[1791] = 10'b0000100001;
mem2[1792] = 10'b0000100010;
mem2[1793] = 10'b0000100010;
mem2[1794] = 10'b0000100010;
mem2[1795] = 10'b0000100010;
mem2[1796] = 10'b0000100010;
mem2[1797] = 10'b0000100010;
mem2[1798] = 10'b0000100010;
mem2[1799] = 10'b0000100010;
mem2[1800] = 10'b0000100010;
mem2[1801] = 10'b0000100010;
mem2[1802] = 10'b0000100010;
mem2[1803] = 10'b0000100010;
mem2[1804] = 10'b0000100010;
mem2[1805] = 10'b0000100010;
mem2[1806] = 10'b0000100010;
mem2[1807] = 10'b0000100010;
mem2[1808] = 10'b0000100010;
mem2[1809] = 10'b0000100010;
mem2[1810] = 10'b0000100010;
mem2[1811] = 10'b0000100010;
mem2[1812] = 10'b0000100010;
mem2[1813] = 10'b0000100010;
mem2[1814] = 10'b0000100010;
mem2[1815] = 10'b0000100010;
mem2[1816] = 10'b0000100010;
mem2[1817] = 10'b0000100010;
mem2[1818] = 10'b0000100011;
mem2[1819] = 10'b0000100011;
mem2[1820] = 10'b0000100011;
mem2[1821] = 10'b0000100011;
mem2[1822] = 10'b0000100011;
mem2[1823] = 10'b0000100011;
mem2[1824] = 10'b0000100011;
mem2[1825] = 10'b0000100011;
mem2[1826] = 10'b0000100011;
mem2[1827] = 10'b0000100011;
mem2[1828] = 10'b0000100011;
mem2[1829] = 10'b0000100011;
mem2[1830] = 10'b0000100011;
mem2[1831] = 10'b0000100011;
mem2[1832] = 10'b0000100011;
mem2[1833] = 10'b0000100011;
mem2[1834] = 10'b0000100011;
mem2[1835] = 10'b0000100011;
mem2[1836] = 10'b0000100011;
mem2[1837] = 10'b0000100011;
mem2[1838] = 10'b0000100011;
mem2[1839] = 10'b0000100011;
mem2[1840] = 10'b0000100011;
mem2[1841] = 10'b0000100011;
mem2[1842] = 10'b0000100011;
mem2[1843] = 10'b0000100011;
mem2[1844] = 10'b0000100011;
mem2[1845] = 10'b0000100100;
mem2[1846] = 10'b0000100100;
mem2[1847] = 10'b0000100100;
mem2[1848] = 10'b0000100100;
mem2[1849] = 10'b0000100100;
mem2[1850] = 10'b0000100100;
mem2[1851] = 10'b0000100100;
mem2[1852] = 10'b0000100100;
mem2[1853] = 10'b0000100100;
mem2[1854] = 10'b0000100100;
mem2[1855] = 10'b0000100100;
mem2[1856] = 10'b0000100100;
mem2[1857] = 10'b0000100100;
mem2[1858] = 10'b0000100100;
mem2[1859] = 10'b0000100100;
mem2[1860] = 10'b0000100100;
mem2[1861] = 10'b0000100100;
mem2[1862] = 10'b0000100100;
mem2[1863] = 10'b0000100100;
mem2[1864] = 10'b0000100100;
mem2[1865] = 10'b0000100100;
mem2[1866] = 10'b0000100100;
mem2[1867] = 10'b0000100100;
mem2[1868] = 10'b0000100100;
mem2[1869] = 10'b0000100100;
mem2[1870] = 10'b0000100101;
mem2[1871] = 10'b0000100101;
mem2[1872] = 10'b0000100101;
mem2[1873] = 10'b0000100101;
mem2[1874] = 10'b0000100101;
mem2[1875] = 10'b0000100101;
mem2[1876] = 10'b0000100101;
mem2[1877] = 10'b0000100101;
mem2[1878] = 10'b0000100101;
mem2[1879] = 10'b0000100101;
mem2[1880] = 10'b0000100101;
mem2[1881] = 10'b0000100101;
mem2[1882] = 10'b0000100101;
mem2[1883] = 10'b0000100101;
mem2[1884] = 10'b0000100101;
mem2[1885] = 10'b0000100101;
mem2[1886] = 10'b0000100101;
mem2[1887] = 10'b0000100101;
mem2[1888] = 10'b0000100101;
mem2[1889] = 10'b0000100101;
mem2[1890] = 10'b0000100101;
mem2[1891] = 10'b0000100101;
mem2[1892] = 10'b0000100101;
mem2[1893] = 10'b0000100101;
mem2[1894] = 10'b0000100101;
mem2[1895] = 10'b0000100101;
mem2[1896] = 10'b0000100110;
mem2[1897] = 10'b0000100110;
mem2[1898] = 10'b0000100110;
mem2[1899] = 10'b0000100110;
mem2[1900] = 10'b0000100110;
mem2[1901] = 10'b0000100110;
mem2[1902] = 10'b0000100110;
mem2[1903] = 10'b0000100110;
mem2[1904] = 10'b0000100110;
mem2[1905] = 10'b0000100110;
mem2[1906] = 10'b0000100110;
mem2[1907] = 10'b0000100110;
mem2[1908] = 10'b0000100110;
mem2[1909] = 10'b0000100110;
mem2[1910] = 10'b0000100110;
mem2[1911] = 10'b0000100110;
mem2[1912] = 10'b0000100110;
mem2[1913] = 10'b0000100110;
mem2[1914] = 10'b0000100110;
mem2[1915] = 10'b0000100110;
mem2[1916] = 10'b0000100110;
mem2[1917] = 10'b0000100110;
mem2[1918] = 10'b0000100110;
mem2[1919] = 10'b0000100110;
mem2[1920] = 10'b0000100110;
mem2[1921] = 10'b0000100111;
mem2[1922] = 10'b0000100111;
mem2[1923] = 10'b0000100111;
mem2[1924] = 10'b0000100111;
mem2[1925] = 10'b0000100111;
mem2[1926] = 10'b0000100111;
mem2[1927] = 10'b0000100111;
mem2[1928] = 10'b0000100111;
mem2[1929] = 10'b0000100111;
mem2[1930] = 10'b0000100111;
mem2[1931] = 10'b0000100111;
mem2[1932] = 10'b0000100111;
mem2[1933] = 10'b0000100111;
mem2[1934] = 10'b0000100111;
mem2[1935] = 10'b0000100111;
mem2[1936] = 10'b0000100111;
mem2[1937] = 10'b0000100111;
mem2[1938] = 10'b0000100111;
mem2[1939] = 10'b0000100111;
mem2[1940] = 10'b0000100111;
mem2[1941] = 10'b0000100111;
mem2[1942] = 10'b0000100111;
mem2[1943] = 10'b0000100111;
mem2[1944] = 10'b0000100111;
mem2[1945] = 10'b0000100111;
mem2[1946] = 10'b0000101000;
mem2[1947] = 10'b0000101000;
mem2[1948] = 10'b0000101000;
mem2[1949] = 10'b0000101000;
mem2[1950] = 10'b0000101000;
mem2[1951] = 10'b0000101000;
mem2[1952] = 10'b0000101000;
mem2[1953] = 10'b0000101000;
mem2[1954] = 10'b0000101000;
mem2[1955] = 10'b0000101000;
mem2[1956] = 10'b0000101000;
mem2[1957] = 10'b0000101000;
mem2[1958] = 10'b0000101000;
mem2[1959] = 10'b0000101000;
mem2[1960] = 10'b0000101000;
mem2[1961] = 10'b0000101000;
mem2[1962] = 10'b0000101000;
mem2[1963] = 10'b0000101000;
mem2[1964] = 10'b0000101000;
mem2[1965] = 10'b0000101000;
mem2[1966] = 10'b0000101000;
mem2[1967] = 10'b0000101000;
mem2[1968] = 10'b0000101000;
mem2[1969] = 10'b0000101000;
mem2[1970] = 10'b0000101001;
mem2[1971] = 10'b0000101001;
mem2[1972] = 10'b0000101001;
mem2[1973] = 10'b0000101001;
mem2[1974] = 10'b0000101001;
mem2[1975] = 10'b0000101001;
mem2[1976] = 10'b0000101001;
mem2[1977] = 10'b0000101001;
mem2[1978] = 10'b0000101001;
mem2[1979] = 10'b0000101001;
mem2[1980] = 10'b0000101001;
mem2[1981] = 10'b0000101001;
mem2[1982] = 10'b0000101001;
mem2[1983] = 10'b0000101001;
mem2[1984] = 10'b0000101001;
mem2[1985] = 10'b0000101001;
mem2[1986] = 10'b0000101001;
mem2[1987] = 10'b0000101001;
mem2[1988] = 10'b0000101001;
mem2[1989] = 10'b0000101001;
mem2[1990] = 10'b0000101001;
mem2[1991] = 10'b0000101001;
mem2[1992] = 10'b0000101001;
mem2[1993] = 10'b0000101001;
mem2[1994] = 10'b0000101010;
mem2[1995] = 10'b0000101010;
mem2[1996] = 10'b0000101010;
mem2[1997] = 10'b0000101010;
mem2[1998] = 10'b0000101010;
mem2[1999] = 10'b0000101010;
mem2[2000] = 10'b0000101010;
mem2[2001] = 10'b0000101010;
mem2[2002] = 10'b0000101010;
mem2[2003] = 10'b0000101010;
mem2[2004] = 10'b0000101010;
mem2[2005] = 10'b0000101010;
mem2[2006] = 10'b0000101010;
mem2[2007] = 10'b0000101010;
mem2[2008] = 10'b0000101010;
mem2[2009] = 10'b0000101010;
mem2[2010] = 10'b0000101010;
mem2[2011] = 10'b0000101010;
mem2[2012] = 10'b0000101010;
mem2[2013] = 10'b0000101010;
mem2[2014] = 10'b0000101010;
mem2[2015] = 10'b0000101010;
mem2[2016] = 10'b0000101010;
mem2[2017] = 10'b0000101010;
mem2[2018] = 10'b0000101011;
mem2[2019] = 10'b0000101011;
mem2[2020] = 10'b0000101011;
mem2[2021] = 10'b0000101011;
mem2[2022] = 10'b0000101011;
mem2[2023] = 10'b0000101011;
mem2[2024] = 10'b0000101011;
mem2[2025] = 10'b0000101011;
mem2[2026] = 10'b0000101011;
mem2[2027] = 10'b0000101011;
mem2[2028] = 10'b0000101011;
mem2[2029] = 10'b0000101011;
mem2[2030] = 10'b0000101011;
mem2[2031] = 10'b0000101011;
mem2[2032] = 10'b0000101011;
mem2[2033] = 10'b0000101011;
mem2[2034] = 10'b0000101011;
mem2[2035] = 10'b0000101011;
mem2[2036] = 10'b0000101011;
mem2[2037] = 10'b0000101011;
mem2[2038] = 10'b0000101011;
mem2[2039] = 10'b0000101011;
mem2[2040] = 10'b0000101011;
mem2[2041] = 10'b0000101011;
mem2[2042] = 10'b0000101100;
mem2[2043] = 10'b0000101100;
mem2[2044] = 10'b0000101100;
mem2[2045] = 10'b0000101100;
mem2[2046] = 10'b0000101100;
mem2[2047] = 10'b0000101100;
mem2[2048] = 10'b0000101100;
mem2[2049] = 10'b0000101100;
mem2[2050] = 10'b0000101100;
mem2[2051] = 10'b0000101100;
mem2[2052] = 10'b0000101100;
mem2[2053] = 10'b0000101100;
mem2[2054] = 10'b0000101100;
mem2[2055] = 10'b0000101100;
mem2[2056] = 10'b0000101100;
mem2[2057] = 10'b0000101100;
mem2[2058] = 10'b0000101100;
mem2[2059] = 10'b0000101100;
mem2[2060] = 10'b0000101100;
mem2[2061] = 10'b0000101100;
mem2[2062] = 10'b0000101100;
mem2[2063] = 10'b0000101100;
mem2[2064] = 10'b0000101100;
mem2[2065] = 10'b0000101101;
mem2[2066] = 10'b0000101101;
mem2[2067] = 10'b0000101101;
mem2[2068] = 10'b0000101101;
mem2[2069] = 10'b0000101101;
mem2[2070] = 10'b0000101101;
mem2[2071] = 10'b0000101101;
mem2[2072] = 10'b0000101101;
mem2[2073] = 10'b0000101101;
mem2[2074] = 10'b0000101101;
mem2[2075] = 10'b0000101101;
mem2[2076] = 10'b0000101101;
mem2[2077] = 10'b0000101101;
mem2[2078] = 10'b0000101101;
mem2[2079] = 10'b0000101101;
mem2[2080] = 10'b0000101101;
mem2[2081] = 10'b0000101101;
mem2[2082] = 10'b0000101101;
mem2[2083] = 10'b0000101101;
mem2[2084] = 10'b0000101101;
mem2[2085] = 10'b0000101101;
mem2[2086] = 10'b0000101101;
mem2[2087] = 10'b0000101101;
mem2[2088] = 10'b0000101101;
mem2[2089] = 10'b0000101110;
mem2[2090] = 10'b0000101110;
mem2[2091] = 10'b0000101110;
mem2[2092] = 10'b0000101110;
mem2[2093] = 10'b0000101110;
mem2[2094] = 10'b0000101110;
mem2[2095] = 10'b0000101110;
mem2[2096] = 10'b0000101110;
mem2[2097] = 10'b0000101110;
mem2[2098] = 10'b0000101110;
mem2[2099] = 10'b0000101110;
mem2[2100] = 10'b0000101110;
mem2[2101] = 10'b0000101110;
mem2[2102] = 10'b0000101110;
mem2[2103] = 10'b0000101110;
mem2[2104] = 10'b0000101110;
mem2[2105] = 10'b0000101110;
mem2[2106] = 10'b0000101110;
mem2[2107] = 10'b0000101110;
mem2[2108] = 10'b0000101110;
mem2[2109] = 10'b0000101110;
mem2[2110] = 10'b0000101110;
mem2[2111] = 10'b0000101111;
mem2[2112] = 10'b0000101111;
mem2[2113] = 10'b0000101111;
mem2[2114] = 10'b0000101111;
mem2[2115] = 10'b0000101111;
mem2[2116] = 10'b0000101111;
mem2[2117] = 10'b0000101111;
mem2[2118] = 10'b0000101111;
mem2[2119] = 10'b0000101111;
mem2[2120] = 10'b0000101111;
mem2[2121] = 10'b0000101111;
mem2[2122] = 10'b0000101111;
mem2[2123] = 10'b0000101111;
mem2[2124] = 10'b0000101111;
mem2[2125] = 10'b0000101111;
mem2[2126] = 10'b0000101111;
mem2[2127] = 10'b0000101111;
mem2[2128] = 10'b0000101111;
mem2[2129] = 10'b0000101111;
mem2[2130] = 10'b0000101111;
mem2[2131] = 10'b0000101111;
mem2[2132] = 10'b0000101111;
mem2[2133] = 10'b0000101111;
mem2[2134] = 10'b0000110000;
mem2[2135] = 10'b0000110000;
mem2[2136] = 10'b0000110000;
mem2[2137] = 10'b0000110000;
mem2[2138] = 10'b0000110000;
mem2[2139] = 10'b0000110000;
mem2[2140] = 10'b0000110000;
mem2[2141] = 10'b0000110000;
mem2[2142] = 10'b0000110000;
mem2[2143] = 10'b0000110000;
mem2[2144] = 10'b0000110000;
mem2[2145] = 10'b0000110000;
mem2[2146] = 10'b0000110000;
mem2[2147] = 10'b0000110000;
mem2[2148] = 10'b0000110000;
mem2[2149] = 10'b0000110000;
mem2[2150] = 10'b0000110000;
mem2[2151] = 10'b0000110000;
mem2[2152] = 10'b0000110000;
mem2[2153] = 10'b0000110000;
mem2[2154] = 10'b0000110000;
mem2[2155] = 10'b0000110000;
mem2[2156] = 10'b0000110000;
mem2[2157] = 10'b0000110001;
mem2[2158] = 10'b0000110001;
mem2[2159] = 10'b0000110001;
mem2[2160] = 10'b0000110001;
mem2[2161] = 10'b0000110001;
mem2[2162] = 10'b0000110001;
mem2[2163] = 10'b0000110001;
mem2[2164] = 10'b0000110001;
mem2[2165] = 10'b0000110001;
mem2[2166] = 10'b0000110001;
mem2[2167] = 10'b0000110001;
mem2[2168] = 10'b0000110001;
mem2[2169] = 10'b0000110001;
mem2[2170] = 10'b0000110001;
mem2[2171] = 10'b0000110001;
mem2[2172] = 10'b0000110001;
mem2[2173] = 10'b0000110001;
mem2[2174] = 10'b0000110001;
mem2[2175] = 10'b0000110001;
mem2[2176] = 10'b0000110001;
mem2[2177] = 10'b0000110001;
mem2[2178] = 10'b0000110001;
mem2[2179] = 10'b0000110010;
mem2[2180] = 10'b0000110010;
mem2[2181] = 10'b0000110010;
mem2[2182] = 10'b0000110010;
mem2[2183] = 10'b0000110010;
mem2[2184] = 10'b0000110010;
mem2[2185] = 10'b0000110010;
mem2[2186] = 10'b0000110010;
mem2[2187] = 10'b0000110010;
mem2[2188] = 10'b0000110010;
mem2[2189] = 10'b0000110010;
mem2[2190] = 10'b0000110010;
mem2[2191] = 10'b0000110010;
mem2[2192] = 10'b0000110010;
mem2[2193] = 10'b0000110010;
mem2[2194] = 10'b0000110010;
mem2[2195] = 10'b0000110010;
mem2[2196] = 10'b0000110010;
mem2[2197] = 10'b0000110010;
mem2[2198] = 10'b0000110010;
mem2[2199] = 10'b0000110010;
mem2[2200] = 10'b0000110010;
mem2[2201] = 10'b0000110011;
mem2[2202] = 10'b0000110011;
mem2[2203] = 10'b0000110011;
mem2[2204] = 10'b0000110011;
mem2[2205] = 10'b0000110011;
mem2[2206] = 10'b0000110011;
mem2[2207] = 10'b0000110011;
mem2[2208] = 10'b0000110011;
mem2[2209] = 10'b0000110011;
mem2[2210] = 10'b0000110011;
mem2[2211] = 10'b0000110011;
mem2[2212] = 10'b0000110011;
mem2[2213] = 10'b0000110011;
mem2[2214] = 10'b0000110011;
mem2[2215] = 10'b0000110011;
mem2[2216] = 10'b0000110011;
mem2[2217] = 10'b0000110011;
mem2[2218] = 10'b0000110011;
mem2[2219] = 10'b0000110011;
mem2[2220] = 10'b0000110011;
mem2[2221] = 10'b0000110011;
mem2[2222] = 10'b0000110011;
mem2[2223] = 10'b0000110100;
mem2[2224] = 10'b0000110100;
mem2[2225] = 10'b0000110100;
mem2[2226] = 10'b0000110100;
mem2[2227] = 10'b0000110100;
mem2[2228] = 10'b0000110100;
mem2[2229] = 10'b0000110100;
mem2[2230] = 10'b0000110100;
mem2[2231] = 10'b0000110100;
mem2[2232] = 10'b0000110100;
mem2[2233] = 10'b0000110100;
mem2[2234] = 10'b0000110100;
mem2[2235] = 10'b0000110100;
mem2[2236] = 10'b0000110100;
mem2[2237] = 10'b0000110100;
mem2[2238] = 10'b0000110100;
mem2[2239] = 10'b0000110100;
mem2[2240] = 10'b0000110100;
mem2[2241] = 10'b0000110100;
mem2[2242] = 10'b0000110100;
mem2[2243] = 10'b0000110100;
mem2[2244] = 10'b0000110101;
mem2[2245] = 10'b0000110101;
mem2[2246] = 10'b0000110101;
mem2[2247] = 10'b0000110101;
mem2[2248] = 10'b0000110101;
mem2[2249] = 10'b0000110101;
mem2[2250] = 10'b0000110101;
mem2[2251] = 10'b0000110101;
mem2[2252] = 10'b0000110101;
mem2[2253] = 10'b0000110101;
mem2[2254] = 10'b0000110101;
mem2[2255] = 10'b0000110101;
mem2[2256] = 10'b0000110101;
mem2[2257] = 10'b0000110101;
mem2[2258] = 10'b0000110101;
mem2[2259] = 10'b0000110101;
mem2[2260] = 10'b0000110101;
mem2[2261] = 10'b0000110101;
mem2[2262] = 10'b0000110101;
mem2[2263] = 10'b0000110101;
mem2[2264] = 10'b0000110101;
mem2[2265] = 10'b0000110101;
mem2[2266] = 10'b0000110110;
mem2[2267] = 10'b0000110110;
mem2[2268] = 10'b0000110110;
mem2[2269] = 10'b0000110110;
mem2[2270] = 10'b0000110110;
mem2[2271] = 10'b0000110110;
mem2[2272] = 10'b0000110110;
mem2[2273] = 10'b0000110110;
mem2[2274] = 10'b0000110110;
mem2[2275] = 10'b0000110110;
mem2[2276] = 10'b0000110110;
mem2[2277] = 10'b0000110110;
mem2[2278] = 10'b0000110110;
mem2[2279] = 10'b0000110110;
mem2[2280] = 10'b0000110110;
mem2[2281] = 10'b0000110110;
mem2[2282] = 10'b0000110110;
mem2[2283] = 10'b0000110110;
mem2[2284] = 10'b0000110110;
mem2[2285] = 10'b0000110110;
mem2[2286] = 10'b0000110110;
mem2[2287] = 10'b0000110111;
mem2[2288] = 10'b0000110111;
mem2[2289] = 10'b0000110111;
mem2[2290] = 10'b0000110111;
mem2[2291] = 10'b0000110111;
mem2[2292] = 10'b0000110111;
mem2[2293] = 10'b0000110111;
mem2[2294] = 10'b0000110111;
mem2[2295] = 10'b0000110111;
mem2[2296] = 10'b0000110111;
mem2[2297] = 10'b0000110111;
mem2[2298] = 10'b0000110111;
mem2[2299] = 10'b0000110111;
mem2[2300] = 10'b0000110111;
mem2[2301] = 10'b0000110111;
mem2[2302] = 10'b0000110111;
mem2[2303] = 10'b0000110111;
mem2[2304] = 10'b0000110111;
mem2[2305] = 10'b0000110111;
mem2[2306] = 10'b0000110111;
mem2[2307] = 10'b0000110111;
mem2[2308] = 10'b0000111000;
mem2[2309] = 10'b0000111000;
mem2[2310] = 10'b0000111000;
mem2[2311] = 10'b0000111000;
mem2[2312] = 10'b0000111000;
mem2[2313] = 10'b0000111000;
mem2[2314] = 10'b0000111000;
mem2[2315] = 10'b0000111000;
mem2[2316] = 10'b0000111000;
mem2[2317] = 10'b0000111000;
mem2[2318] = 10'b0000111000;
mem2[2319] = 10'b0000111000;
mem2[2320] = 10'b0000111000;
mem2[2321] = 10'b0000111000;
mem2[2322] = 10'b0000111000;
mem2[2323] = 10'b0000111000;
mem2[2324] = 10'b0000111000;
mem2[2325] = 10'b0000111000;
mem2[2326] = 10'b0000111000;
mem2[2327] = 10'b0000111000;
mem2[2328] = 10'b0000111000;
mem2[2329] = 10'b0000111001;
mem2[2330] = 10'b0000111001;
mem2[2331] = 10'b0000111001;
mem2[2332] = 10'b0000111001;
mem2[2333] = 10'b0000111001;
mem2[2334] = 10'b0000111001;
mem2[2335] = 10'b0000111001;
mem2[2336] = 10'b0000111001;
mem2[2337] = 10'b0000111001;
mem2[2338] = 10'b0000111001;
mem2[2339] = 10'b0000111001;
mem2[2340] = 10'b0000111001;
mem2[2341] = 10'b0000111001;
mem2[2342] = 10'b0000111001;
mem2[2343] = 10'b0000111001;
mem2[2344] = 10'b0000111001;
mem2[2345] = 10'b0000111001;
mem2[2346] = 10'b0000111001;
mem2[2347] = 10'b0000111001;
mem2[2348] = 10'b0000111001;
mem2[2349] = 10'b0000111001;
mem2[2350] = 10'b0000111010;
mem2[2351] = 10'b0000111010;
mem2[2352] = 10'b0000111010;
mem2[2353] = 10'b0000111010;
mem2[2354] = 10'b0000111010;
mem2[2355] = 10'b0000111010;
mem2[2356] = 10'b0000111010;
mem2[2357] = 10'b0000111010;
mem2[2358] = 10'b0000111010;
mem2[2359] = 10'b0000111010;
mem2[2360] = 10'b0000111010;
mem2[2361] = 10'b0000111010;
mem2[2362] = 10'b0000111010;
mem2[2363] = 10'b0000111010;
mem2[2364] = 10'b0000111010;
mem2[2365] = 10'b0000111010;
mem2[2366] = 10'b0000111010;
mem2[2367] = 10'b0000111010;
mem2[2368] = 10'b0000111010;
mem2[2369] = 10'b0000111010;
mem2[2370] = 10'b0000111010;
mem2[2371] = 10'b0000111011;
mem2[2372] = 10'b0000111011;
mem2[2373] = 10'b0000111011;
mem2[2374] = 10'b0000111011;
mem2[2375] = 10'b0000111011;
mem2[2376] = 10'b0000111011;
mem2[2377] = 10'b0000111011;
mem2[2378] = 10'b0000111011;
mem2[2379] = 10'b0000111011;
mem2[2380] = 10'b0000111011;
mem2[2381] = 10'b0000111011;
mem2[2382] = 10'b0000111011;
mem2[2383] = 10'b0000111011;
mem2[2384] = 10'b0000111011;
mem2[2385] = 10'b0000111011;
mem2[2386] = 10'b0000111011;
mem2[2387] = 10'b0000111011;
mem2[2388] = 10'b0000111011;
mem2[2389] = 10'b0000111011;
mem2[2390] = 10'b0000111011;
mem2[2391] = 10'b0000111100;
mem2[2392] = 10'b0000111100;
mem2[2393] = 10'b0000111100;
mem2[2394] = 10'b0000111100;
mem2[2395] = 10'b0000111100;
mem2[2396] = 10'b0000111100;
mem2[2397] = 10'b0000111100;
mem2[2398] = 10'b0000111100;
mem2[2399] = 10'b0000111100;
mem2[2400] = 10'b0000111100;
mem2[2401] = 10'b0000111100;
mem2[2402] = 10'b0000111100;
mem2[2403] = 10'b0000111100;
mem2[2404] = 10'b0000111100;
mem2[2405] = 10'b0000111100;
mem2[2406] = 10'b0000111100;
mem2[2407] = 10'b0000111100;
mem2[2408] = 10'b0000111100;
mem2[2409] = 10'b0000111100;
mem2[2410] = 10'b0000111100;
mem2[2411] = 10'b0000111101;
mem2[2412] = 10'b0000111101;
mem2[2413] = 10'b0000111101;
mem2[2414] = 10'b0000111101;
mem2[2415] = 10'b0000111101;
mem2[2416] = 10'b0000111101;
mem2[2417] = 10'b0000111101;
mem2[2418] = 10'b0000111101;
mem2[2419] = 10'b0000111101;
mem2[2420] = 10'b0000111101;
mem2[2421] = 10'b0000111101;
mem2[2422] = 10'b0000111101;
mem2[2423] = 10'b0000111101;
mem2[2424] = 10'b0000111101;
mem2[2425] = 10'b0000111101;
mem2[2426] = 10'b0000111101;
mem2[2427] = 10'b0000111101;
mem2[2428] = 10'b0000111101;
mem2[2429] = 10'b0000111101;
mem2[2430] = 10'b0000111101;
mem2[2431] = 10'b0000111110;
mem2[2432] = 10'b0000111110;
mem2[2433] = 10'b0000111110;
mem2[2434] = 10'b0000111110;
mem2[2435] = 10'b0000111110;
mem2[2436] = 10'b0000111110;
mem2[2437] = 10'b0000111110;
mem2[2438] = 10'b0000111110;
mem2[2439] = 10'b0000111110;
mem2[2440] = 10'b0000111110;
mem2[2441] = 10'b0000111110;
mem2[2442] = 10'b0000111110;
mem2[2443] = 10'b0000111110;
mem2[2444] = 10'b0000111110;
mem2[2445] = 10'b0000111110;
mem2[2446] = 10'b0000111110;
mem2[2447] = 10'b0000111110;
mem2[2448] = 10'b0000111110;
mem2[2449] = 10'b0000111110;
mem2[2450] = 10'b0000111110;
mem2[2451] = 10'b0000111111;
mem2[2452] = 10'b0000111111;
mem2[2453] = 10'b0000111111;
mem2[2454] = 10'b0000111111;
mem2[2455] = 10'b0000111111;
mem2[2456] = 10'b0000111111;
mem2[2457] = 10'b0000111111;
mem2[2458] = 10'b0000111111;
mem2[2459] = 10'b0000111111;
mem2[2460] = 10'b0000111111;
mem2[2461] = 10'b0000111111;
mem2[2462] = 10'b0000111111;
mem2[2463] = 10'b0000111111;
mem2[2464] = 10'b0000111111;
mem2[2465] = 10'b0000111111;
mem2[2466] = 10'b0000111111;
mem2[2467] = 10'b0000111111;
mem2[2468] = 10'b0000111111;
mem2[2469] = 10'b0000111111;
mem2[2470] = 10'b0000111111;
mem2[2471] = 10'b0001000000;
mem2[2472] = 10'b0001000000;
mem2[2473] = 10'b0001000000;
mem2[2474] = 10'b0001000000;
mem2[2475] = 10'b0001000000;
mem2[2476] = 10'b0001000000;
mem2[2477] = 10'b0001000000;
mem2[2478] = 10'b0001000000;
mem2[2479] = 10'b0001000000;
mem2[2480] = 10'b0001000000;
mem2[2481] = 10'b0001000000;
mem2[2482] = 10'b0001000000;
mem2[2483] = 10'b0001000000;
mem2[2484] = 10'b0001000000;
mem2[2485] = 10'b0001000000;
mem2[2486] = 10'b0001000000;
mem2[2487] = 10'b0001000000;
mem2[2488] = 10'b0001000000;
mem2[2489] = 10'b0001000000;
mem2[2490] = 10'b0001000000;
mem2[2491] = 10'b0001000001;
mem2[2492] = 10'b0001000001;
mem2[2493] = 10'b0001000001;
mem2[2494] = 10'b0001000001;
mem2[2495] = 10'b0001000001;
mem2[2496] = 10'b0001000001;
mem2[2497] = 10'b0001000001;
mem2[2498] = 10'b0001000001;
mem2[2499] = 10'b0001000001;
mem2[2500] = 10'b0001000001;
mem2[2501] = 10'b0001000001;
mem2[2502] = 10'b0001000001;
mem2[2503] = 10'b0001000001;
mem2[2504] = 10'b0001000001;
mem2[2505] = 10'b0001000001;
mem2[2506] = 10'b0001000001;
mem2[2507] = 10'b0001000001;
mem2[2508] = 10'b0001000001;
mem2[2509] = 10'b0001000001;
mem2[2510] = 10'b0001000010;
mem2[2511] = 10'b0001000010;
mem2[2512] = 10'b0001000010;
mem2[2513] = 10'b0001000010;
mem2[2514] = 10'b0001000010;
mem2[2515] = 10'b0001000010;
mem2[2516] = 10'b0001000010;
mem2[2517] = 10'b0001000010;
mem2[2518] = 10'b0001000010;
mem2[2519] = 10'b0001000010;
mem2[2520] = 10'b0001000010;
mem2[2521] = 10'b0001000010;
mem2[2522] = 10'b0001000010;
mem2[2523] = 10'b0001000010;
mem2[2524] = 10'b0001000010;
mem2[2525] = 10'b0001000010;
mem2[2526] = 10'b0001000010;
mem2[2527] = 10'b0001000010;
mem2[2528] = 10'b0001000010;
mem2[2529] = 10'b0001000010;
mem2[2530] = 10'b0001000011;
mem2[2531] = 10'b0001000011;
mem2[2532] = 10'b0001000011;
mem2[2533] = 10'b0001000011;
mem2[2534] = 10'b0001000011;
mem2[2535] = 10'b0001000011;
mem2[2536] = 10'b0001000011;
mem2[2537] = 10'b0001000011;
mem2[2538] = 10'b0001000011;
mem2[2539] = 10'b0001000011;
mem2[2540] = 10'b0001000011;
mem2[2541] = 10'b0001000011;
mem2[2542] = 10'b0001000011;
mem2[2543] = 10'b0001000011;
mem2[2544] = 10'b0001000011;
mem2[2545] = 10'b0001000011;
mem2[2546] = 10'b0001000011;
mem2[2547] = 10'b0001000011;
mem2[2548] = 10'b0001000011;
mem2[2549] = 10'b0001000100;
mem2[2550] = 10'b0001000100;
mem2[2551] = 10'b0001000100;
mem2[2552] = 10'b0001000100;
mem2[2553] = 10'b0001000100;
mem2[2554] = 10'b0001000100;
mem2[2555] = 10'b0001000100;
mem2[2556] = 10'b0001000100;
mem2[2557] = 10'b0001000100;
mem2[2558] = 10'b0001000100;
mem2[2559] = 10'b0001000100;
mem2[2560] = 10'b0001000100;
mem2[2561] = 10'b0001000100;
mem2[2562] = 10'b0001000100;
mem2[2563] = 10'b0001000100;
mem2[2564] = 10'b0001000100;
mem2[2565] = 10'b0001000100;
mem2[2566] = 10'b0001000100;
mem2[2567] = 10'b0001000100;
mem2[2568] = 10'b0001000101;
mem2[2569] = 10'b0001000101;
mem2[2570] = 10'b0001000101;
mem2[2571] = 10'b0001000101;
mem2[2572] = 10'b0001000101;
mem2[2573] = 10'b0001000101;
mem2[2574] = 10'b0001000101;
mem2[2575] = 10'b0001000101;
mem2[2576] = 10'b0001000101;
mem2[2577] = 10'b0001000101;
mem2[2578] = 10'b0001000101;
mem2[2579] = 10'b0001000101;
mem2[2580] = 10'b0001000101;
mem2[2581] = 10'b0001000101;
mem2[2582] = 10'b0001000101;
mem2[2583] = 10'b0001000101;
mem2[2584] = 10'b0001000101;
mem2[2585] = 10'b0001000101;
mem2[2586] = 10'b0001000101;
mem2[2587] = 10'b0001000110;
mem2[2588] = 10'b0001000110;
mem2[2589] = 10'b0001000110;
mem2[2590] = 10'b0001000110;
mem2[2591] = 10'b0001000110;
mem2[2592] = 10'b0001000110;
mem2[2593] = 10'b0001000110;
mem2[2594] = 10'b0001000110;
mem2[2595] = 10'b0001000110;
mem2[2596] = 10'b0001000110;
mem2[2597] = 10'b0001000110;
mem2[2598] = 10'b0001000110;
mem2[2599] = 10'b0001000110;
mem2[2600] = 10'b0001000110;
mem2[2601] = 10'b0001000110;
mem2[2602] = 10'b0001000110;
mem2[2603] = 10'b0001000110;
mem2[2604] = 10'b0001000110;
mem2[2605] = 10'b0001000110;
mem2[2606] = 10'b0001000111;
mem2[2607] = 10'b0001000111;
mem2[2608] = 10'b0001000111;
mem2[2609] = 10'b0001000111;
mem2[2610] = 10'b0001000111;
mem2[2611] = 10'b0001000111;
mem2[2612] = 10'b0001000111;
mem2[2613] = 10'b0001000111;
mem2[2614] = 10'b0001000111;
mem2[2615] = 10'b0001000111;
mem2[2616] = 10'b0001000111;
mem2[2617] = 10'b0001000111;
mem2[2618] = 10'b0001000111;
mem2[2619] = 10'b0001000111;
mem2[2620] = 10'b0001000111;
mem2[2621] = 10'b0001000111;
mem2[2622] = 10'b0001000111;
mem2[2623] = 10'b0001000111;
mem2[2624] = 10'b0001001000;
mem2[2625] = 10'b0001001000;
mem2[2626] = 10'b0001001000;
mem2[2627] = 10'b0001001000;
mem2[2628] = 10'b0001001000;
mem2[2629] = 10'b0001001000;
mem2[2630] = 10'b0001001000;
mem2[2631] = 10'b0001001000;
mem2[2632] = 10'b0001001000;
mem2[2633] = 10'b0001001000;
mem2[2634] = 10'b0001001000;
mem2[2635] = 10'b0001001000;
mem2[2636] = 10'b0001001000;
mem2[2637] = 10'b0001001000;
mem2[2638] = 10'b0001001000;
mem2[2639] = 10'b0001001000;
mem2[2640] = 10'b0001001000;
mem2[2641] = 10'b0001001000;
mem2[2642] = 10'b0001001000;
mem2[2643] = 10'b0001001001;
mem2[2644] = 10'b0001001001;
mem2[2645] = 10'b0001001001;
mem2[2646] = 10'b0001001001;
mem2[2647] = 10'b0001001001;
mem2[2648] = 10'b0001001001;
mem2[2649] = 10'b0001001001;
mem2[2650] = 10'b0001001001;
mem2[2651] = 10'b0001001001;
mem2[2652] = 10'b0001001001;
mem2[2653] = 10'b0001001001;
mem2[2654] = 10'b0001001001;
mem2[2655] = 10'b0001001001;
mem2[2656] = 10'b0001001001;
mem2[2657] = 10'b0001001001;
mem2[2658] = 10'b0001001001;
mem2[2659] = 10'b0001001001;
mem2[2660] = 10'b0001001001;
mem2[2661] = 10'b0001001001;
mem2[2662] = 10'b0001001010;
mem2[2663] = 10'b0001001010;
mem2[2664] = 10'b0001001010;
mem2[2665] = 10'b0001001010;
mem2[2666] = 10'b0001001010;
mem2[2667] = 10'b0001001010;
mem2[2668] = 10'b0001001010;
mem2[2669] = 10'b0001001010;
mem2[2670] = 10'b0001001010;
mem2[2671] = 10'b0001001010;
mem2[2672] = 10'b0001001010;
mem2[2673] = 10'b0001001010;
mem2[2674] = 10'b0001001010;
mem2[2675] = 10'b0001001010;
mem2[2676] = 10'b0001001010;
mem2[2677] = 10'b0001001010;
mem2[2678] = 10'b0001001010;
mem2[2679] = 10'b0001001010;
mem2[2680] = 10'b0001001011;
mem2[2681] = 10'b0001001011;
mem2[2682] = 10'b0001001011;
mem2[2683] = 10'b0001001011;
mem2[2684] = 10'b0001001011;
mem2[2685] = 10'b0001001011;
mem2[2686] = 10'b0001001011;
mem2[2687] = 10'b0001001011;
mem2[2688] = 10'b0001001011;
mem2[2689] = 10'b0001001011;
mem2[2690] = 10'b0001001011;
mem2[2691] = 10'b0001001011;
mem2[2692] = 10'b0001001011;
mem2[2693] = 10'b0001001011;
mem2[2694] = 10'b0001001011;
mem2[2695] = 10'b0001001011;
mem2[2696] = 10'b0001001011;
mem2[2697] = 10'b0001001011;
mem2[2698] = 10'b0001001100;
mem2[2699] = 10'b0001001100;
mem2[2700] = 10'b0001001100;
mem2[2701] = 10'b0001001100;
mem2[2702] = 10'b0001001100;
mem2[2703] = 10'b0001001100;
mem2[2704] = 10'b0001001100;
mem2[2705] = 10'b0001001100;
mem2[2706] = 10'b0001001100;
mem2[2707] = 10'b0001001100;
mem2[2708] = 10'b0001001100;
mem2[2709] = 10'b0001001100;
mem2[2710] = 10'b0001001100;
mem2[2711] = 10'b0001001100;
mem2[2712] = 10'b0001001100;
mem2[2713] = 10'b0001001100;
mem2[2714] = 10'b0001001100;
mem2[2715] = 10'b0001001100;
mem2[2716] = 10'b0001001101;
mem2[2717] = 10'b0001001101;
mem2[2718] = 10'b0001001101;
mem2[2719] = 10'b0001001101;
mem2[2720] = 10'b0001001101;
mem2[2721] = 10'b0001001101;
mem2[2722] = 10'b0001001101;
mem2[2723] = 10'b0001001101;
mem2[2724] = 10'b0001001101;
mem2[2725] = 10'b0001001101;
mem2[2726] = 10'b0001001101;
mem2[2727] = 10'b0001001101;
mem2[2728] = 10'b0001001101;
mem2[2729] = 10'b0001001101;
mem2[2730] = 10'b0001001101;
mem2[2731] = 10'b0001001101;
mem2[2732] = 10'b0001001101;
mem2[2733] = 10'b0001001101;
mem2[2734] = 10'b0001001110;
mem2[2735] = 10'b0001001110;
mem2[2736] = 10'b0001001110;
mem2[2737] = 10'b0001001110;
mem2[2738] = 10'b0001001110;
mem2[2739] = 10'b0001001110;
mem2[2740] = 10'b0001001110;
mem2[2741] = 10'b0001001110;
mem2[2742] = 10'b0001001110;
mem2[2743] = 10'b0001001110;
mem2[2744] = 10'b0001001110;
mem2[2745] = 10'b0001001110;
mem2[2746] = 10'b0001001110;
mem2[2747] = 10'b0001001110;
mem2[2748] = 10'b0001001110;
mem2[2749] = 10'b0001001110;
mem2[2750] = 10'b0001001110;
mem2[2751] = 10'b0001001110;
mem2[2752] = 10'b0001001111;
mem2[2753] = 10'b0001001111;
mem2[2754] = 10'b0001001111;
mem2[2755] = 10'b0001001111;
mem2[2756] = 10'b0001001111;
mem2[2757] = 10'b0001001111;
mem2[2758] = 10'b0001001111;
mem2[2759] = 10'b0001001111;
mem2[2760] = 10'b0001001111;
mem2[2761] = 10'b0001001111;
mem2[2762] = 10'b0001001111;
mem2[2763] = 10'b0001001111;
mem2[2764] = 10'b0001001111;
mem2[2765] = 10'b0001001111;
mem2[2766] = 10'b0001001111;
mem2[2767] = 10'b0001001111;
mem2[2768] = 10'b0001001111;
mem2[2769] = 10'b0001001111;
mem2[2770] = 10'b0001010000;
mem2[2771] = 10'b0001010000;
mem2[2772] = 10'b0001010000;
mem2[2773] = 10'b0001010000;
mem2[2774] = 10'b0001010000;
mem2[2775] = 10'b0001010000;
mem2[2776] = 10'b0001010000;
mem2[2777] = 10'b0001010000;
mem2[2778] = 10'b0001010000;
mem2[2779] = 10'b0001010000;
mem2[2780] = 10'b0001010000;
mem2[2781] = 10'b0001010000;
mem2[2782] = 10'b0001010000;
mem2[2783] = 10'b0001010000;
mem2[2784] = 10'b0001010000;
mem2[2785] = 10'b0001010000;
mem2[2786] = 10'b0001010000;
mem2[2787] = 10'b0001010000;
mem2[2788] = 10'b0001010001;
mem2[2789] = 10'b0001010001;
mem2[2790] = 10'b0001010001;
mem2[2791] = 10'b0001010001;
mem2[2792] = 10'b0001010001;
mem2[2793] = 10'b0001010001;
mem2[2794] = 10'b0001010001;
mem2[2795] = 10'b0001010001;
mem2[2796] = 10'b0001010001;
mem2[2797] = 10'b0001010001;
mem2[2798] = 10'b0001010001;
mem2[2799] = 10'b0001010001;
mem2[2800] = 10'b0001010001;
mem2[2801] = 10'b0001010001;
mem2[2802] = 10'b0001010001;
mem2[2803] = 10'b0001010001;
mem2[2804] = 10'b0001010001;
mem2[2805] = 10'b0001010001;
mem2[2806] = 10'b0001010010;
mem2[2807] = 10'b0001010010;
mem2[2808] = 10'b0001010010;
mem2[2809] = 10'b0001010010;
mem2[2810] = 10'b0001010010;
mem2[2811] = 10'b0001010010;
mem2[2812] = 10'b0001010010;
mem2[2813] = 10'b0001010010;
mem2[2814] = 10'b0001010010;
mem2[2815] = 10'b0001010010;
mem2[2816] = 10'b0001010010;
mem2[2817] = 10'b0001010010;
mem2[2818] = 10'b0001010010;
mem2[2819] = 10'b0001010010;
mem2[2820] = 10'b0001010010;
mem2[2821] = 10'b0001010010;
mem2[2822] = 10'b0001010010;
mem2[2823] = 10'b0001010011;
mem2[2824] = 10'b0001010011;
mem2[2825] = 10'b0001010011;
mem2[2826] = 10'b0001010011;
mem2[2827] = 10'b0001010011;
mem2[2828] = 10'b0001010011;
mem2[2829] = 10'b0001010011;
mem2[2830] = 10'b0001010011;
mem2[2831] = 10'b0001010011;
mem2[2832] = 10'b0001010011;
mem2[2833] = 10'b0001010011;
mem2[2834] = 10'b0001010011;
mem2[2835] = 10'b0001010011;
mem2[2836] = 10'b0001010011;
mem2[2837] = 10'b0001010011;
mem2[2838] = 10'b0001010011;
mem2[2839] = 10'b0001010011;
mem2[2840] = 10'b0001010011;
mem2[2841] = 10'b0001010100;
mem2[2842] = 10'b0001010100;
mem2[2843] = 10'b0001010100;
mem2[2844] = 10'b0001010100;
mem2[2845] = 10'b0001010100;
mem2[2846] = 10'b0001010100;
mem2[2847] = 10'b0001010100;
mem2[2848] = 10'b0001010100;
mem2[2849] = 10'b0001010100;
mem2[2850] = 10'b0001010100;
mem2[2851] = 10'b0001010100;
mem2[2852] = 10'b0001010100;
mem2[2853] = 10'b0001010100;
mem2[2854] = 10'b0001010100;
mem2[2855] = 10'b0001010100;
mem2[2856] = 10'b0001010100;
mem2[2857] = 10'b0001010100;
mem2[2858] = 10'b0001010101;
mem2[2859] = 10'b0001010101;
mem2[2860] = 10'b0001010101;
mem2[2861] = 10'b0001010101;
mem2[2862] = 10'b0001010101;
mem2[2863] = 10'b0001010101;
mem2[2864] = 10'b0001010101;
mem2[2865] = 10'b0001010101;
mem2[2866] = 10'b0001010101;
mem2[2867] = 10'b0001010101;
mem2[2868] = 10'b0001010101;
mem2[2869] = 10'b0001010101;
mem2[2870] = 10'b0001010101;
mem2[2871] = 10'b0001010101;
mem2[2872] = 10'b0001010101;
mem2[2873] = 10'b0001010101;
mem2[2874] = 10'b0001010101;
mem2[2875] = 10'b0001010110;
mem2[2876] = 10'b0001010110;
mem2[2877] = 10'b0001010110;
mem2[2878] = 10'b0001010110;
mem2[2879] = 10'b0001010110;
mem2[2880] = 10'b0001010110;
mem2[2881] = 10'b0001010110;
mem2[2882] = 10'b0001010110;
mem2[2883] = 10'b0001010110;
mem2[2884] = 10'b0001010110;
mem2[2885] = 10'b0001010110;
mem2[2886] = 10'b0001010110;
mem2[2887] = 10'b0001010110;
mem2[2888] = 10'b0001010110;
mem2[2889] = 10'b0001010110;
mem2[2890] = 10'b0001010110;
mem2[2891] = 10'b0001010110;
mem2[2892] = 10'b0001010111;
mem2[2893] = 10'b0001010111;
mem2[2894] = 10'b0001010111;
mem2[2895] = 10'b0001010111;
mem2[2896] = 10'b0001010111;
mem2[2897] = 10'b0001010111;
mem2[2898] = 10'b0001010111;
mem2[2899] = 10'b0001010111;
mem2[2900] = 10'b0001010111;
mem2[2901] = 10'b0001010111;
mem2[2902] = 10'b0001010111;
mem2[2903] = 10'b0001010111;
mem2[2904] = 10'b0001010111;
mem2[2905] = 10'b0001010111;
mem2[2906] = 10'b0001010111;
mem2[2907] = 10'b0001010111;
mem2[2908] = 10'b0001010111;
mem2[2909] = 10'b0001011000;
mem2[2910] = 10'b0001011000;
mem2[2911] = 10'b0001011000;
mem2[2912] = 10'b0001011000;
mem2[2913] = 10'b0001011000;
mem2[2914] = 10'b0001011000;
mem2[2915] = 10'b0001011000;
mem2[2916] = 10'b0001011000;
mem2[2917] = 10'b0001011000;
mem2[2918] = 10'b0001011000;
mem2[2919] = 10'b0001011000;
mem2[2920] = 10'b0001011000;
mem2[2921] = 10'b0001011000;
mem2[2922] = 10'b0001011000;
mem2[2923] = 10'b0001011000;
mem2[2924] = 10'b0001011000;
mem2[2925] = 10'b0001011000;
mem2[2926] = 10'b0001011001;
mem2[2927] = 10'b0001011001;
mem2[2928] = 10'b0001011001;
mem2[2929] = 10'b0001011001;
mem2[2930] = 10'b0001011001;
mem2[2931] = 10'b0001011001;
mem2[2932] = 10'b0001011001;
mem2[2933] = 10'b0001011001;
mem2[2934] = 10'b0001011001;
mem2[2935] = 10'b0001011001;
mem2[2936] = 10'b0001011001;
mem2[2937] = 10'b0001011001;
mem2[2938] = 10'b0001011001;
mem2[2939] = 10'b0001011001;
mem2[2940] = 10'b0001011001;
mem2[2941] = 10'b0001011001;
mem2[2942] = 10'b0001011001;
mem2[2943] = 10'b0001011010;
mem2[2944] = 10'b0001011010;
mem2[2945] = 10'b0001011010;
mem2[2946] = 10'b0001011010;
mem2[2947] = 10'b0001011010;
mem2[2948] = 10'b0001011010;
mem2[2949] = 10'b0001011010;
mem2[2950] = 10'b0001011010;
mem2[2951] = 10'b0001011010;
mem2[2952] = 10'b0001011010;
mem2[2953] = 10'b0001011010;
mem2[2954] = 10'b0001011010;
mem2[2955] = 10'b0001011010;
mem2[2956] = 10'b0001011010;
mem2[2957] = 10'b0001011010;
mem2[2958] = 10'b0001011010;
mem2[2959] = 10'b0001011010;
mem2[2960] = 10'b0001011011;
mem2[2961] = 10'b0001011011;
mem2[2962] = 10'b0001011011;
mem2[2963] = 10'b0001011011;
mem2[2964] = 10'b0001011011;
mem2[2965] = 10'b0001011011;
mem2[2966] = 10'b0001011011;
mem2[2967] = 10'b0001011011;
mem2[2968] = 10'b0001011011;
mem2[2969] = 10'b0001011011;
mem2[2970] = 10'b0001011011;
mem2[2971] = 10'b0001011011;
mem2[2972] = 10'b0001011011;
mem2[2973] = 10'b0001011011;
mem2[2974] = 10'b0001011011;
mem2[2975] = 10'b0001011011;
mem2[2976] = 10'b0001011011;
mem2[2977] = 10'b0001011100;
mem2[2978] = 10'b0001011100;
mem2[2979] = 10'b0001011100;
mem2[2980] = 10'b0001011100;
mem2[2981] = 10'b0001011100;
mem2[2982] = 10'b0001011100;
mem2[2983] = 10'b0001011100;
mem2[2984] = 10'b0001011100;
mem2[2985] = 10'b0001011100;
mem2[2986] = 10'b0001011100;
mem2[2987] = 10'b0001011100;
mem2[2988] = 10'b0001011100;
mem2[2989] = 10'b0001011100;
mem2[2990] = 10'b0001011100;
mem2[2991] = 10'b0001011100;
mem2[2992] = 10'b0001011100;
mem2[2993] = 10'b0001011100;
mem2[2994] = 10'b0001011101;
mem2[2995] = 10'b0001011101;
mem2[2996] = 10'b0001011101;
mem2[2997] = 10'b0001011101;
mem2[2998] = 10'b0001011101;
mem2[2999] = 10'b0001011101;
mem2[3000] = 10'b0001011101;
mem2[3001] = 10'b0001011101;
mem2[3002] = 10'b0001011101;
mem2[3003] = 10'b0001011101;
mem2[3004] = 10'b0001011101;
mem2[3005] = 10'b0001011101;
mem2[3006] = 10'b0001011101;
mem2[3007] = 10'b0001011101;
mem2[3008] = 10'b0001011101;
mem2[3009] = 10'b0001011101;
mem2[3010] = 10'b0001011110;
mem2[3011] = 10'b0001011110;
mem2[3012] = 10'b0001011110;
mem2[3013] = 10'b0001011110;
mem2[3014] = 10'b0001011110;
mem2[3015] = 10'b0001011110;
mem2[3016] = 10'b0001011110;
mem2[3017] = 10'b0001011110;
mem2[3018] = 10'b0001011110;
mem2[3019] = 10'b0001011110;
mem2[3020] = 10'b0001011110;
mem2[3021] = 10'b0001011110;
mem2[3022] = 10'b0001011110;
mem2[3023] = 10'b0001011110;
mem2[3024] = 10'b0001011110;
mem2[3025] = 10'b0001011110;
mem2[3026] = 10'b0001011110;
mem2[3027] = 10'b0001011111;
mem2[3028] = 10'b0001011111;
mem2[3029] = 10'b0001011111;
mem2[3030] = 10'b0001011111;
mem2[3031] = 10'b0001011111;
mem2[3032] = 10'b0001011111;
mem2[3033] = 10'b0001011111;
mem2[3034] = 10'b0001011111;
mem2[3035] = 10'b0001011111;
mem2[3036] = 10'b0001011111;
mem2[3037] = 10'b0001011111;
mem2[3038] = 10'b0001011111;
mem2[3039] = 10'b0001011111;
mem2[3040] = 10'b0001011111;
mem2[3041] = 10'b0001011111;
mem2[3042] = 10'b0001011111;
mem2[3043] = 10'b0001100000;
mem2[3044] = 10'b0001100000;
mem2[3045] = 10'b0001100000;
mem2[3046] = 10'b0001100000;
mem2[3047] = 10'b0001100000;
mem2[3048] = 10'b0001100000;
mem2[3049] = 10'b0001100000;
mem2[3050] = 10'b0001100000;
mem2[3051] = 10'b0001100000;
mem2[3052] = 10'b0001100000;
mem2[3053] = 10'b0001100000;
mem2[3054] = 10'b0001100000;
mem2[3055] = 10'b0001100000;
mem2[3056] = 10'b0001100000;
mem2[3057] = 10'b0001100000;
mem2[3058] = 10'b0001100000;
mem2[3059] = 10'b0001100001;
mem2[3060] = 10'b0001100001;
mem2[3061] = 10'b0001100001;
mem2[3062] = 10'b0001100001;
mem2[3063] = 10'b0001100001;
mem2[3064] = 10'b0001100001;
mem2[3065] = 10'b0001100001;
mem2[3066] = 10'b0001100001;
mem2[3067] = 10'b0001100001;
mem2[3068] = 10'b0001100001;
mem2[3069] = 10'b0001100001;
mem2[3070] = 10'b0001100001;
mem2[3071] = 10'b0001100001;
mem2[3072] = 10'b0001100001;
mem2[3073] = 10'b0001100001;
mem2[3074] = 10'b0001100001;
mem2[3075] = 10'b0001100001;
mem2[3076] = 10'b0001100010;
mem2[3077] = 10'b0001100010;
mem2[3078] = 10'b0001100010;
mem2[3079] = 10'b0001100010;
mem2[3080] = 10'b0001100010;
mem2[3081] = 10'b0001100010;
mem2[3082] = 10'b0001100010;
mem2[3083] = 10'b0001100010;
mem2[3084] = 10'b0001100010;
mem2[3085] = 10'b0001100010;
mem2[3086] = 10'b0001100010;
mem2[3087] = 10'b0001100010;
mem2[3088] = 10'b0001100010;
mem2[3089] = 10'b0001100010;
mem2[3090] = 10'b0001100010;
mem2[3091] = 10'b0001100010;
mem2[3092] = 10'b0001100011;
mem2[3093] = 10'b0001100011;
mem2[3094] = 10'b0001100011;
mem2[3095] = 10'b0001100011;
mem2[3096] = 10'b0001100011;
mem2[3097] = 10'b0001100011;
mem2[3098] = 10'b0001100011;
mem2[3099] = 10'b0001100011;
mem2[3100] = 10'b0001100011;
mem2[3101] = 10'b0001100011;
mem2[3102] = 10'b0001100011;
mem2[3103] = 10'b0001100011;
mem2[3104] = 10'b0001100011;
mem2[3105] = 10'b0001100011;
mem2[3106] = 10'b0001100011;
mem2[3107] = 10'b0001100011;
mem2[3108] = 10'b0001100100;
mem2[3109] = 10'b0001100100;
mem2[3110] = 10'b0001100100;
mem2[3111] = 10'b0001100100;
mem2[3112] = 10'b0001100100;
mem2[3113] = 10'b0001100100;
mem2[3114] = 10'b0001100100;
mem2[3115] = 10'b0001100100;
mem2[3116] = 10'b0001100100;
mem2[3117] = 10'b0001100100;
mem2[3118] = 10'b0001100100;
mem2[3119] = 10'b0001100100;
mem2[3120] = 10'b0001100100;
mem2[3121] = 10'b0001100100;
mem2[3122] = 10'b0001100100;
mem2[3123] = 10'b0001100100;
mem2[3124] = 10'b0001100101;
mem2[3125] = 10'b0001100101;
mem2[3126] = 10'b0001100101;
mem2[3127] = 10'b0001100101;
mem2[3128] = 10'b0001100101;
mem2[3129] = 10'b0001100101;
mem2[3130] = 10'b0001100101;
mem2[3131] = 10'b0001100101;
mem2[3132] = 10'b0001100101;
mem2[3133] = 10'b0001100101;
mem2[3134] = 10'b0001100101;
mem2[3135] = 10'b0001100101;
mem2[3136] = 10'b0001100101;
mem2[3137] = 10'b0001100101;
mem2[3138] = 10'b0001100101;
mem2[3139] = 10'b0001100101;
mem2[3140] = 10'b0001100110;
mem2[3141] = 10'b0001100110;
mem2[3142] = 10'b0001100110;
mem2[3143] = 10'b0001100110;
mem2[3144] = 10'b0001100110;
mem2[3145] = 10'b0001100110;
mem2[3146] = 10'b0001100110;
mem2[3147] = 10'b0001100110;
mem2[3148] = 10'b0001100110;
mem2[3149] = 10'b0001100110;
mem2[3150] = 10'b0001100110;
mem2[3151] = 10'b0001100110;
mem2[3152] = 10'b0001100110;
mem2[3153] = 10'b0001100110;
mem2[3154] = 10'b0001100110;
mem2[3155] = 10'b0001100110;
mem2[3156] = 10'b0001100111;
mem2[3157] = 10'b0001100111;
mem2[3158] = 10'b0001100111;
mem2[3159] = 10'b0001100111;
mem2[3160] = 10'b0001100111;
mem2[3161] = 10'b0001100111;
mem2[3162] = 10'b0001100111;
mem2[3163] = 10'b0001100111;
mem2[3164] = 10'b0001100111;
mem2[3165] = 10'b0001100111;
mem2[3166] = 10'b0001100111;
mem2[3167] = 10'b0001100111;
mem2[3168] = 10'b0001100111;
mem2[3169] = 10'b0001100111;
mem2[3170] = 10'b0001100111;
mem2[3171] = 10'b0001100111;
mem2[3172] = 10'b0001101000;
mem2[3173] = 10'b0001101000;
mem2[3174] = 10'b0001101000;
mem2[3175] = 10'b0001101000;
mem2[3176] = 10'b0001101000;
mem2[3177] = 10'b0001101000;
mem2[3178] = 10'b0001101000;
mem2[3179] = 10'b0001101000;
mem2[3180] = 10'b0001101000;
mem2[3181] = 10'b0001101000;
mem2[3182] = 10'b0001101000;
mem2[3183] = 10'b0001101000;
mem2[3184] = 10'b0001101000;
mem2[3185] = 10'b0001101000;
mem2[3186] = 10'b0001101000;
mem2[3187] = 10'b0001101000;
mem2[3188] = 10'b0001101001;
mem2[3189] = 10'b0001101001;
mem2[3190] = 10'b0001101001;
mem2[3191] = 10'b0001101001;
mem2[3192] = 10'b0001101001;
mem2[3193] = 10'b0001101001;
mem2[3194] = 10'b0001101001;
mem2[3195] = 10'b0001101001;
mem2[3196] = 10'b0001101001;
mem2[3197] = 10'b0001101001;
mem2[3198] = 10'b0001101001;
mem2[3199] = 10'b0001101001;
mem2[3200] = 10'b0001101001;
mem2[3201] = 10'b0001101001;
mem2[3202] = 10'b0001101001;
mem2[3203] = 10'b0001101010;
mem2[3204] = 10'b0001101010;
mem2[3205] = 10'b0001101010;
mem2[3206] = 10'b0001101010;
mem2[3207] = 10'b0001101010;
mem2[3208] = 10'b0001101010;
mem2[3209] = 10'b0001101010;
mem2[3210] = 10'b0001101010;
mem2[3211] = 10'b0001101010;
mem2[3212] = 10'b0001101010;
mem2[3213] = 10'b0001101010;
mem2[3214] = 10'b0001101010;
mem2[3215] = 10'b0001101010;
mem2[3216] = 10'b0001101010;
mem2[3217] = 10'b0001101010;
mem2[3218] = 10'b0001101010;
mem2[3219] = 10'b0001101011;
mem2[3220] = 10'b0001101011;
mem2[3221] = 10'b0001101011;
mem2[3222] = 10'b0001101011;
mem2[3223] = 10'b0001101011;
mem2[3224] = 10'b0001101011;
mem2[3225] = 10'b0001101011;
mem2[3226] = 10'b0001101011;
mem2[3227] = 10'b0001101011;
mem2[3228] = 10'b0001101011;
mem2[3229] = 10'b0001101011;
mem2[3230] = 10'b0001101011;
mem2[3231] = 10'b0001101011;
mem2[3232] = 10'b0001101011;
mem2[3233] = 10'b0001101011;
mem2[3234] = 10'b0001101100;
mem2[3235] = 10'b0001101100;
mem2[3236] = 10'b0001101100;
mem2[3237] = 10'b0001101100;
mem2[3238] = 10'b0001101100;
mem2[3239] = 10'b0001101100;
mem2[3240] = 10'b0001101100;
mem2[3241] = 10'b0001101100;
mem2[3242] = 10'b0001101100;
mem2[3243] = 10'b0001101100;
mem2[3244] = 10'b0001101100;
mem2[3245] = 10'b0001101100;
mem2[3246] = 10'b0001101100;
mem2[3247] = 10'b0001101100;
mem2[3248] = 10'b0001101100;
mem2[3249] = 10'b0001101100;
mem2[3250] = 10'b0001101101;
mem2[3251] = 10'b0001101101;
mem2[3252] = 10'b0001101101;
mem2[3253] = 10'b0001101101;
mem2[3254] = 10'b0001101101;
mem2[3255] = 10'b0001101101;
mem2[3256] = 10'b0001101101;
mem2[3257] = 10'b0001101101;
mem2[3258] = 10'b0001101101;
mem2[3259] = 10'b0001101101;
mem2[3260] = 10'b0001101101;
mem2[3261] = 10'b0001101101;
mem2[3262] = 10'b0001101101;
mem2[3263] = 10'b0001101101;
mem2[3264] = 10'b0001101101;
mem2[3265] = 10'b0001101110;
mem2[3266] = 10'b0001101110;
mem2[3267] = 10'b0001101110;
mem2[3268] = 10'b0001101110;
mem2[3269] = 10'b0001101110;
mem2[3270] = 10'b0001101110;
mem2[3271] = 10'b0001101110;
mem2[3272] = 10'b0001101110;
mem2[3273] = 10'b0001101110;
mem2[3274] = 10'b0001101110;
mem2[3275] = 10'b0001101110;
mem2[3276] = 10'b0001101110;
mem2[3277] = 10'b0001101110;
mem2[3278] = 10'b0001101110;
mem2[3279] = 10'b0001101110;
mem2[3280] = 10'b0001101110;
mem2[3281] = 10'b0001101111;
mem2[3282] = 10'b0001101111;
mem2[3283] = 10'b0001101111;
mem2[3284] = 10'b0001101111;
mem2[3285] = 10'b0001101111;
mem2[3286] = 10'b0001101111;
mem2[3287] = 10'b0001101111;
mem2[3288] = 10'b0001101111;
mem2[3289] = 10'b0001101111;
mem2[3290] = 10'b0001101111;
mem2[3291] = 10'b0001101111;
mem2[3292] = 10'b0001101111;
mem2[3293] = 10'b0001101111;
mem2[3294] = 10'b0001101111;
mem2[3295] = 10'b0001101111;
mem2[3296] = 10'b0001110000;
mem2[3297] = 10'b0001110000;
mem2[3298] = 10'b0001110000;
mem2[3299] = 10'b0001110000;
mem2[3300] = 10'b0001110000;
mem2[3301] = 10'b0001110000;
mem2[3302] = 10'b0001110000;
mem2[3303] = 10'b0001110000;
mem2[3304] = 10'b0001110000;
mem2[3305] = 10'b0001110000;
mem2[3306] = 10'b0001110000;
mem2[3307] = 10'b0001110000;
mem2[3308] = 10'b0001110000;
mem2[3309] = 10'b0001110000;
mem2[3310] = 10'b0001110000;
mem2[3311] = 10'b0001110001;
mem2[3312] = 10'b0001110001;
mem2[3313] = 10'b0001110001;
mem2[3314] = 10'b0001110001;
mem2[3315] = 10'b0001110001;
mem2[3316] = 10'b0001110001;
mem2[3317] = 10'b0001110001;
mem2[3318] = 10'b0001110001;
mem2[3319] = 10'b0001110001;
mem2[3320] = 10'b0001110001;
mem2[3321] = 10'b0001110001;
mem2[3322] = 10'b0001110001;
mem2[3323] = 10'b0001110001;
mem2[3324] = 10'b0001110001;
mem2[3325] = 10'b0001110001;
mem2[3326] = 10'b0001110001;
mem2[3327] = 10'b0001110010;
mem2[3328] = 10'b0001110010;
mem2[3329] = 10'b0001110010;
mem2[3330] = 10'b0001110010;
mem2[3331] = 10'b0001110010;
mem2[3332] = 10'b0001110010;
mem2[3333] = 10'b0001110010;
mem2[3334] = 10'b0001110010;
mem2[3335] = 10'b0001110010;
mem2[3336] = 10'b0001110010;
mem2[3337] = 10'b0001110010;
mem2[3338] = 10'b0001110010;
mem2[3339] = 10'b0001110010;
mem2[3340] = 10'b0001110010;
mem2[3341] = 10'b0001110010;
mem2[3342] = 10'b0001110011;
mem2[3343] = 10'b0001110011;
mem2[3344] = 10'b0001110011;
mem2[3345] = 10'b0001110011;
mem2[3346] = 10'b0001110011;
mem2[3347] = 10'b0001110011;
mem2[3348] = 10'b0001110011;
mem2[3349] = 10'b0001110011;
mem2[3350] = 10'b0001110011;
mem2[3351] = 10'b0001110011;
mem2[3352] = 10'b0001110011;
mem2[3353] = 10'b0001110011;
mem2[3354] = 10'b0001110011;
mem2[3355] = 10'b0001110011;
mem2[3356] = 10'b0001110011;
mem2[3357] = 10'b0001110100;
mem2[3358] = 10'b0001110100;
mem2[3359] = 10'b0001110100;
mem2[3360] = 10'b0001110100;
mem2[3361] = 10'b0001110100;
mem2[3362] = 10'b0001110100;
mem2[3363] = 10'b0001110100;
mem2[3364] = 10'b0001110100;
mem2[3365] = 10'b0001110100;
mem2[3366] = 10'b0001110100;
mem2[3367] = 10'b0001110100;
mem2[3368] = 10'b0001110100;
mem2[3369] = 10'b0001110100;
mem2[3370] = 10'b0001110100;
mem2[3371] = 10'b0001110100;
mem2[3372] = 10'b0001110101;
mem2[3373] = 10'b0001110101;
mem2[3374] = 10'b0001110101;
mem2[3375] = 10'b0001110101;
mem2[3376] = 10'b0001110101;
mem2[3377] = 10'b0001110101;
mem2[3378] = 10'b0001110101;
mem2[3379] = 10'b0001110101;
mem2[3380] = 10'b0001110101;
mem2[3381] = 10'b0001110101;
mem2[3382] = 10'b0001110101;
mem2[3383] = 10'b0001110101;
mem2[3384] = 10'b0001110101;
mem2[3385] = 10'b0001110101;
mem2[3386] = 10'b0001110101;
mem2[3387] = 10'b0001110110;
mem2[3388] = 10'b0001110110;
mem2[3389] = 10'b0001110110;
mem2[3390] = 10'b0001110110;
mem2[3391] = 10'b0001110110;
mem2[3392] = 10'b0001110110;
mem2[3393] = 10'b0001110110;
mem2[3394] = 10'b0001110110;
mem2[3395] = 10'b0001110110;
mem2[3396] = 10'b0001110110;
mem2[3397] = 10'b0001110110;
mem2[3398] = 10'b0001110110;
mem2[3399] = 10'b0001110110;
mem2[3400] = 10'b0001110110;
mem2[3401] = 10'b0001110110;
mem2[3402] = 10'b0001110111;
mem2[3403] = 10'b0001110111;
mem2[3404] = 10'b0001110111;
mem2[3405] = 10'b0001110111;
mem2[3406] = 10'b0001110111;
mem2[3407] = 10'b0001110111;
mem2[3408] = 10'b0001110111;
mem2[3409] = 10'b0001110111;
mem2[3410] = 10'b0001110111;
mem2[3411] = 10'b0001110111;
mem2[3412] = 10'b0001110111;
mem2[3413] = 10'b0001110111;
mem2[3414] = 10'b0001110111;
mem2[3415] = 10'b0001110111;
mem2[3416] = 10'b0001110111;
mem2[3417] = 10'b0001111000;
mem2[3418] = 10'b0001111000;
mem2[3419] = 10'b0001111000;
mem2[3420] = 10'b0001111000;
mem2[3421] = 10'b0001111000;
mem2[3422] = 10'b0001111000;
mem2[3423] = 10'b0001111000;
mem2[3424] = 10'b0001111000;
mem2[3425] = 10'b0001111000;
mem2[3426] = 10'b0001111000;
mem2[3427] = 10'b0001111000;
mem2[3428] = 10'b0001111000;
mem2[3429] = 10'b0001111000;
mem2[3430] = 10'b0001111000;
mem2[3431] = 10'b0001111001;
mem2[3432] = 10'b0001111001;
mem2[3433] = 10'b0001111001;
mem2[3434] = 10'b0001111001;
mem2[3435] = 10'b0001111001;
mem2[3436] = 10'b0001111001;
mem2[3437] = 10'b0001111001;
mem2[3438] = 10'b0001111001;
mem2[3439] = 10'b0001111001;
mem2[3440] = 10'b0001111001;
mem2[3441] = 10'b0001111001;
mem2[3442] = 10'b0001111001;
mem2[3443] = 10'b0001111001;
mem2[3444] = 10'b0001111001;
mem2[3445] = 10'b0001111001;
mem2[3446] = 10'b0001111010;
mem2[3447] = 10'b0001111010;
mem2[3448] = 10'b0001111010;
mem2[3449] = 10'b0001111010;
mem2[3450] = 10'b0001111010;
mem2[3451] = 10'b0001111010;
mem2[3452] = 10'b0001111010;
mem2[3453] = 10'b0001111010;
mem2[3454] = 10'b0001111010;
mem2[3455] = 10'b0001111010;
mem2[3456] = 10'b0001111010;
mem2[3457] = 10'b0001111010;
mem2[3458] = 10'b0001111010;
mem2[3459] = 10'b0001111010;
mem2[3460] = 10'b0001111010;
mem2[3461] = 10'b0001111011;
mem2[3462] = 10'b0001111011;
mem2[3463] = 10'b0001111011;
mem2[3464] = 10'b0001111011;
mem2[3465] = 10'b0001111011;
mem2[3466] = 10'b0001111011;
mem2[3467] = 10'b0001111011;
mem2[3468] = 10'b0001111011;
mem2[3469] = 10'b0001111011;
mem2[3470] = 10'b0001111011;
mem2[3471] = 10'b0001111011;
mem2[3472] = 10'b0001111011;
mem2[3473] = 10'b0001111011;
mem2[3474] = 10'b0001111011;
mem2[3475] = 10'b0001111011;
mem2[3476] = 10'b0001111100;
mem2[3477] = 10'b0001111100;
mem2[3478] = 10'b0001111100;
mem2[3479] = 10'b0001111100;
mem2[3480] = 10'b0001111100;
mem2[3481] = 10'b0001111100;
mem2[3482] = 10'b0001111100;
mem2[3483] = 10'b0001111100;
mem2[3484] = 10'b0001111100;
mem2[3485] = 10'b0001111100;
mem2[3486] = 10'b0001111100;
mem2[3487] = 10'b0001111100;
mem2[3488] = 10'b0001111100;
mem2[3489] = 10'b0001111100;
mem2[3490] = 10'b0001111101;
mem2[3491] = 10'b0001111101;
mem2[3492] = 10'b0001111101;
mem2[3493] = 10'b0001111101;
mem2[3494] = 10'b0001111101;
mem2[3495] = 10'b0001111101;
mem2[3496] = 10'b0001111101;
mem2[3497] = 10'b0001111101;
mem2[3498] = 10'b0001111101;
mem2[3499] = 10'b0001111101;
mem2[3500] = 10'b0001111101;
mem2[3501] = 10'b0001111101;
mem2[3502] = 10'b0001111101;
mem2[3503] = 10'b0001111101;
mem2[3504] = 10'b0001111101;
mem2[3505] = 10'b0001111110;
mem2[3506] = 10'b0001111110;
mem2[3507] = 10'b0001111110;
mem2[3508] = 10'b0001111110;
mem2[3509] = 10'b0001111110;
mem2[3510] = 10'b0001111110;
mem2[3511] = 10'b0001111110;
mem2[3512] = 10'b0001111110;
mem2[3513] = 10'b0001111110;
mem2[3514] = 10'b0001111110;
mem2[3515] = 10'b0001111110;
mem2[3516] = 10'b0001111110;
mem2[3517] = 10'b0001111110;
mem2[3518] = 10'b0001111110;
mem2[3519] = 10'b0001111111;
mem2[3520] = 10'b0001111111;
mem2[3521] = 10'b0001111111;
mem2[3522] = 10'b0001111111;
mem2[3523] = 10'b0001111111;
mem2[3524] = 10'b0001111111;
mem2[3525] = 10'b0001111111;
mem2[3526] = 10'b0001111111;
mem2[3527] = 10'b0001111111;
mem2[3528] = 10'b0001111111;
mem2[3529] = 10'b0001111111;
mem2[3530] = 10'b0001111111;
mem2[3531] = 10'b0001111111;
mem2[3532] = 10'b0001111111;
mem2[3533] = 10'b0001111111;
mem2[3534] = 10'b0010000000;
mem2[3535] = 10'b0010000000;
mem2[3536] = 10'b0010000000;
mem2[3537] = 10'b0010000000;
mem2[3538] = 10'b0010000000;
mem2[3539] = 10'b0010000000;
mem2[3540] = 10'b0010000000;
mem2[3541] = 10'b0010000000;
mem2[3542] = 10'b0010000000;
mem2[3543] = 10'b0010000000;
mem2[3544] = 10'b0010000000;
mem2[3545] = 10'b0010000000;
mem2[3546] = 10'b0010000000;
mem2[3547] = 10'b0010000000;
mem2[3548] = 10'b0010000001;
mem2[3549] = 10'b0010000001;
mem2[3550] = 10'b0010000001;
mem2[3551] = 10'b0010000001;
mem2[3552] = 10'b0010000001;
mem2[3553] = 10'b0010000001;
mem2[3554] = 10'b0010000001;
mem2[3555] = 10'b0010000001;
mem2[3556] = 10'b0010000001;
mem2[3557] = 10'b0010000001;
mem2[3558] = 10'b0010000001;
mem2[3559] = 10'b0010000001;
mem2[3560] = 10'b0010000001;
mem2[3561] = 10'b0010000001;
mem2[3562] = 10'b0010000001;
mem2[3563] = 10'b0010000010;
mem2[3564] = 10'b0010000010;
mem2[3565] = 10'b0010000010;
mem2[3566] = 10'b0010000010;
mem2[3567] = 10'b0010000010;
mem2[3568] = 10'b0010000010;
mem2[3569] = 10'b0010000010;
mem2[3570] = 10'b0010000010;
mem2[3571] = 10'b0010000010;
mem2[3572] = 10'b0010000010;
mem2[3573] = 10'b0010000010;
mem2[3574] = 10'b0010000010;
mem2[3575] = 10'b0010000010;
mem2[3576] = 10'b0010000010;
mem2[3577] = 10'b0010000011;
mem2[3578] = 10'b0010000011;
mem2[3579] = 10'b0010000011;
mem2[3580] = 10'b0010000011;
mem2[3581] = 10'b0010000011;
mem2[3582] = 10'b0010000011;
mem2[3583] = 10'b0010000011;
mem2[3584] = 10'b0010000011;
mem2[3585] = 10'b0010000011;
mem2[3586] = 10'b0010000011;
mem2[3587] = 10'b0010000011;
mem2[3588] = 10'b0010000011;
mem2[3589] = 10'b0010000011;
mem2[3590] = 10'b0010000011;
mem2[3591] = 10'b0010000100;
mem2[3592] = 10'b0010000100;
mem2[3593] = 10'b0010000100;
mem2[3594] = 10'b0010000100;
mem2[3595] = 10'b0010000100;
mem2[3596] = 10'b0010000100;
mem2[3597] = 10'b0010000100;
mem2[3598] = 10'b0010000100;
mem2[3599] = 10'b0010000100;
mem2[3600] = 10'b0010000100;
mem2[3601] = 10'b0010000100;
mem2[3602] = 10'b0010000100;
mem2[3603] = 10'b0010000100;
mem2[3604] = 10'b0010000100;
mem2[3605] = 10'b0010000101;
mem2[3606] = 10'b0010000101;
mem2[3607] = 10'b0010000101;
mem2[3608] = 10'b0010000101;
mem2[3609] = 10'b0010000101;
mem2[3610] = 10'b0010000101;
mem2[3611] = 10'b0010000101;
mem2[3612] = 10'b0010000101;
mem2[3613] = 10'b0010000101;
mem2[3614] = 10'b0010000101;
mem2[3615] = 10'b0010000101;
mem2[3616] = 10'b0010000101;
mem2[3617] = 10'b0010000101;
mem2[3618] = 10'b0010000101;
mem2[3619] = 10'b0010000101;
mem2[3620] = 10'b0010000110;
mem2[3621] = 10'b0010000110;
mem2[3622] = 10'b0010000110;
mem2[3623] = 10'b0010000110;
mem2[3624] = 10'b0010000110;
mem2[3625] = 10'b0010000110;
mem2[3626] = 10'b0010000110;
mem2[3627] = 10'b0010000110;
mem2[3628] = 10'b0010000110;
mem2[3629] = 10'b0010000110;
mem2[3630] = 10'b0010000110;
mem2[3631] = 10'b0010000110;
mem2[3632] = 10'b0010000110;
mem2[3633] = 10'b0010000110;
mem2[3634] = 10'b0010000111;
mem2[3635] = 10'b0010000111;
mem2[3636] = 10'b0010000111;
mem2[3637] = 10'b0010000111;
mem2[3638] = 10'b0010000111;
mem2[3639] = 10'b0010000111;
mem2[3640] = 10'b0010000111;
mem2[3641] = 10'b0010000111;
mem2[3642] = 10'b0010000111;
mem2[3643] = 10'b0010000111;
mem2[3644] = 10'b0010000111;
mem2[3645] = 10'b0010000111;
mem2[3646] = 10'b0010000111;
mem2[3647] = 10'b0010000111;
mem2[3648] = 10'b0010001000;
mem2[3649] = 10'b0010001000;
mem2[3650] = 10'b0010001000;
mem2[3651] = 10'b0010001000;
mem2[3652] = 10'b0010001000;
mem2[3653] = 10'b0010001000;
mem2[3654] = 10'b0010001000;
mem2[3655] = 10'b0010001000;
mem2[3656] = 10'b0010001000;
mem2[3657] = 10'b0010001000;
mem2[3658] = 10'b0010001000;
mem2[3659] = 10'b0010001000;
mem2[3660] = 10'b0010001000;
mem2[3661] = 10'b0010001000;
mem2[3662] = 10'b0010001001;
mem2[3663] = 10'b0010001001;
mem2[3664] = 10'b0010001001;
mem2[3665] = 10'b0010001001;
mem2[3666] = 10'b0010001001;
mem2[3667] = 10'b0010001001;
mem2[3668] = 10'b0010001001;
mem2[3669] = 10'b0010001001;
mem2[3670] = 10'b0010001001;
mem2[3671] = 10'b0010001001;
mem2[3672] = 10'b0010001001;
mem2[3673] = 10'b0010001001;
mem2[3674] = 10'b0010001001;
mem2[3675] = 10'b0010001001;
mem2[3676] = 10'b0010001010;
mem2[3677] = 10'b0010001010;
mem2[3678] = 10'b0010001010;
mem2[3679] = 10'b0010001010;
mem2[3680] = 10'b0010001010;
mem2[3681] = 10'b0010001010;
mem2[3682] = 10'b0010001010;
mem2[3683] = 10'b0010001010;
mem2[3684] = 10'b0010001010;
mem2[3685] = 10'b0010001010;
mem2[3686] = 10'b0010001010;
mem2[3687] = 10'b0010001010;
mem2[3688] = 10'b0010001010;
mem2[3689] = 10'b0010001010;
mem2[3690] = 10'b0010001011;
mem2[3691] = 10'b0010001011;
mem2[3692] = 10'b0010001011;
mem2[3693] = 10'b0010001011;
mem2[3694] = 10'b0010001011;
mem2[3695] = 10'b0010001011;
mem2[3696] = 10'b0010001011;
mem2[3697] = 10'b0010001011;
mem2[3698] = 10'b0010001011;
mem2[3699] = 10'b0010001011;
mem2[3700] = 10'b0010001011;
mem2[3701] = 10'b0010001011;
mem2[3702] = 10'b0010001011;
mem2[3703] = 10'b0010001011;
mem2[3704] = 10'b0010001100;
mem2[3705] = 10'b0010001100;
mem2[3706] = 10'b0010001100;
mem2[3707] = 10'b0010001100;
mem2[3708] = 10'b0010001100;
mem2[3709] = 10'b0010001100;
mem2[3710] = 10'b0010001100;
mem2[3711] = 10'b0010001100;
mem2[3712] = 10'b0010001100;
mem2[3713] = 10'b0010001100;
mem2[3714] = 10'b0010001100;
mem2[3715] = 10'b0010001100;
mem2[3716] = 10'b0010001100;
mem2[3717] = 10'b0010001100;
mem2[3718] = 10'b0010001101;
mem2[3719] = 10'b0010001101;
mem2[3720] = 10'b0010001101;
mem2[3721] = 10'b0010001101;
mem2[3722] = 10'b0010001101;
mem2[3723] = 10'b0010001101;
mem2[3724] = 10'b0010001101;
mem2[3725] = 10'b0010001101;
mem2[3726] = 10'b0010001101;
mem2[3727] = 10'b0010001101;
mem2[3728] = 10'b0010001101;
mem2[3729] = 10'b0010001101;
mem2[3730] = 10'b0010001101;
mem2[3731] = 10'b0010001110;
mem2[3732] = 10'b0010001110;
mem2[3733] = 10'b0010001110;
mem2[3734] = 10'b0010001110;
mem2[3735] = 10'b0010001110;
mem2[3736] = 10'b0010001110;
mem2[3737] = 10'b0010001110;
mem2[3738] = 10'b0010001110;
mem2[3739] = 10'b0010001110;
mem2[3740] = 10'b0010001110;
mem2[3741] = 10'b0010001110;
mem2[3742] = 10'b0010001110;
mem2[3743] = 10'b0010001110;
mem2[3744] = 10'b0010001110;
mem2[3745] = 10'b0010001111;
mem2[3746] = 10'b0010001111;
mem2[3747] = 10'b0010001111;
mem2[3748] = 10'b0010001111;
mem2[3749] = 10'b0010001111;
mem2[3750] = 10'b0010001111;
mem2[3751] = 10'b0010001111;
mem2[3752] = 10'b0010001111;
mem2[3753] = 10'b0010001111;
mem2[3754] = 10'b0010001111;
mem2[3755] = 10'b0010001111;
mem2[3756] = 10'b0010001111;
mem2[3757] = 10'b0010001111;
mem2[3758] = 10'b0010001111;
mem2[3759] = 10'b0010010000;
mem2[3760] = 10'b0010010000;
mem2[3761] = 10'b0010010000;
mem2[3762] = 10'b0010010000;
mem2[3763] = 10'b0010010000;
mem2[3764] = 10'b0010010000;
mem2[3765] = 10'b0010010000;
mem2[3766] = 10'b0010010000;
mem2[3767] = 10'b0010010000;
mem2[3768] = 10'b0010010000;
mem2[3769] = 10'b0010010000;
mem2[3770] = 10'b0010010000;
mem2[3771] = 10'b0010010000;
mem2[3772] = 10'b0010010000;
mem2[3773] = 10'b0010010001;
mem2[3774] = 10'b0010010001;
mem2[3775] = 10'b0010010001;
mem2[3776] = 10'b0010010001;
mem2[3777] = 10'b0010010001;
mem2[3778] = 10'b0010010001;
mem2[3779] = 10'b0010010001;
mem2[3780] = 10'b0010010001;
mem2[3781] = 10'b0010010001;
mem2[3782] = 10'b0010010001;
mem2[3783] = 10'b0010010001;
mem2[3784] = 10'b0010010001;
mem2[3785] = 10'b0010010001;
mem2[3786] = 10'b0010010010;
mem2[3787] = 10'b0010010010;
mem2[3788] = 10'b0010010010;
mem2[3789] = 10'b0010010010;
mem2[3790] = 10'b0010010010;
mem2[3791] = 10'b0010010010;
mem2[3792] = 10'b0010010010;
mem2[3793] = 10'b0010010010;
mem2[3794] = 10'b0010010010;
mem2[3795] = 10'b0010010010;
mem2[3796] = 10'b0010010010;
mem2[3797] = 10'b0010010010;
mem2[3798] = 10'b0010010010;
mem2[3799] = 10'b0010010010;
mem2[3800] = 10'b0010010011;
mem2[3801] = 10'b0010010011;
mem2[3802] = 10'b0010010011;
mem2[3803] = 10'b0010010011;
mem2[3804] = 10'b0010010011;
mem2[3805] = 10'b0010010011;
mem2[3806] = 10'b0010010011;
mem2[3807] = 10'b0010010011;
mem2[3808] = 10'b0010010011;
mem2[3809] = 10'b0010010011;
mem2[3810] = 10'b0010010011;
mem2[3811] = 10'b0010010011;
mem2[3812] = 10'b0010010011;
mem2[3813] = 10'b0010010011;
mem2[3814] = 10'b0010010100;
mem2[3815] = 10'b0010010100;
mem2[3816] = 10'b0010010100;
mem2[3817] = 10'b0010010100;
mem2[3818] = 10'b0010010100;
mem2[3819] = 10'b0010010100;
mem2[3820] = 10'b0010010100;
mem2[3821] = 10'b0010010100;
mem2[3822] = 10'b0010010100;
mem2[3823] = 10'b0010010100;
mem2[3824] = 10'b0010010100;
mem2[3825] = 10'b0010010100;
mem2[3826] = 10'b0010010100;
mem2[3827] = 10'b0010010101;
mem2[3828] = 10'b0010010101;
mem2[3829] = 10'b0010010101;
mem2[3830] = 10'b0010010101;
mem2[3831] = 10'b0010010101;
mem2[3832] = 10'b0010010101;
mem2[3833] = 10'b0010010101;
mem2[3834] = 10'b0010010101;
mem2[3835] = 10'b0010010101;
mem2[3836] = 10'b0010010101;
mem2[3837] = 10'b0010010101;
mem2[3838] = 10'b0010010101;
mem2[3839] = 10'b0010010101;
mem2[3840] = 10'b0010010101;
mem2[3841] = 10'b0010010110;
mem2[3842] = 10'b0010010110;
mem2[3843] = 10'b0010010110;
mem2[3844] = 10'b0010010110;
mem2[3845] = 10'b0010010110;
mem2[3846] = 10'b0010010110;
mem2[3847] = 10'b0010010110;
mem2[3848] = 10'b0010010110;
mem2[3849] = 10'b0010010110;
mem2[3850] = 10'b0010010110;
mem2[3851] = 10'b0010010110;
mem2[3852] = 10'b0010010110;
mem2[3853] = 10'b0010010110;
mem2[3854] = 10'b0010010111;
mem2[3855] = 10'b0010010111;
mem2[3856] = 10'b0010010111;
mem2[3857] = 10'b0010010111;
mem2[3858] = 10'b0010010111;
mem2[3859] = 10'b0010010111;
mem2[3860] = 10'b0010010111;
mem2[3861] = 10'b0010010111;
mem2[3862] = 10'b0010010111;
mem2[3863] = 10'b0010010111;
mem2[3864] = 10'b0010010111;
mem2[3865] = 10'b0010010111;
mem2[3866] = 10'b0010010111;
mem2[3867] = 10'b0010010111;
mem2[3868] = 10'b0010011000;
mem2[3869] = 10'b0010011000;
mem2[3870] = 10'b0010011000;
mem2[3871] = 10'b0010011000;
mem2[3872] = 10'b0010011000;
mem2[3873] = 10'b0010011000;
mem2[3874] = 10'b0010011000;
mem2[3875] = 10'b0010011000;
mem2[3876] = 10'b0010011000;
mem2[3877] = 10'b0010011000;
mem2[3878] = 10'b0010011000;
mem2[3879] = 10'b0010011000;
mem2[3880] = 10'b0010011000;
mem2[3881] = 10'b0010011001;
mem2[3882] = 10'b0010011001;
mem2[3883] = 10'b0010011001;
mem2[3884] = 10'b0010011001;
mem2[3885] = 10'b0010011001;
mem2[3886] = 10'b0010011001;
mem2[3887] = 10'b0010011001;
mem2[3888] = 10'b0010011001;
mem2[3889] = 10'b0010011001;
mem2[3890] = 10'b0010011001;
mem2[3891] = 10'b0010011001;
mem2[3892] = 10'b0010011001;
mem2[3893] = 10'b0010011001;
mem2[3894] = 10'b0010011010;
mem2[3895] = 10'b0010011010;
mem2[3896] = 10'b0010011010;
mem2[3897] = 10'b0010011010;
mem2[3898] = 10'b0010011010;
mem2[3899] = 10'b0010011010;
mem2[3900] = 10'b0010011010;
mem2[3901] = 10'b0010011010;
mem2[3902] = 10'b0010011010;
mem2[3903] = 10'b0010011010;
mem2[3904] = 10'b0010011010;
mem2[3905] = 10'b0010011010;
mem2[3906] = 10'b0010011010;
mem2[3907] = 10'b0010011010;
mem2[3908] = 10'b0010011011;
mem2[3909] = 10'b0010011011;
mem2[3910] = 10'b0010011011;
mem2[3911] = 10'b0010011011;
mem2[3912] = 10'b0010011011;
mem2[3913] = 10'b0010011011;
mem2[3914] = 10'b0010011011;
mem2[3915] = 10'b0010011011;
mem2[3916] = 10'b0010011011;
mem2[3917] = 10'b0010011011;
mem2[3918] = 10'b0010011011;
mem2[3919] = 10'b0010011011;
mem2[3920] = 10'b0010011011;
mem2[3921] = 10'b0010011100;
mem2[3922] = 10'b0010011100;
mem2[3923] = 10'b0010011100;
mem2[3924] = 10'b0010011100;
mem2[3925] = 10'b0010011100;
mem2[3926] = 10'b0010011100;
mem2[3927] = 10'b0010011100;
mem2[3928] = 10'b0010011100;
mem2[3929] = 10'b0010011100;
mem2[3930] = 10'b0010011100;
mem2[3931] = 10'b0010011100;
mem2[3932] = 10'b0010011100;
mem2[3933] = 10'b0010011100;
mem2[3934] = 10'b0010011101;
mem2[3935] = 10'b0010011101;
mem2[3936] = 10'b0010011101;
mem2[3937] = 10'b0010011101;
mem2[3938] = 10'b0010011101;
mem2[3939] = 10'b0010011101;
mem2[3940] = 10'b0010011101;
mem2[3941] = 10'b0010011101;
mem2[3942] = 10'b0010011101;
mem2[3943] = 10'b0010011101;
mem2[3944] = 10'b0010011101;
mem2[3945] = 10'b0010011101;
mem2[3946] = 10'b0010011101;
mem2[3947] = 10'b0010011101;
mem2[3948] = 10'b0010011110;
mem2[3949] = 10'b0010011110;
mem2[3950] = 10'b0010011110;
mem2[3951] = 10'b0010011110;
mem2[3952] = 10'b0010011110;
mem2[3953] = 10'b0010011110;
mem2[3954] = 10'b0010011110;
mem2[3955] = 10'b0010011110;
mem2[3956] = 10'b0010011110;
mem2[3957] = 10'b0010011110;
mem2[3958] = 10'b0010011110;
mem2[3959] = 10'b0010011110;
mem2[3960] = 10'b0010011110;
mem2[3961] = 10'b0010011111;
mem2[3962] = 10'b0010011111;
mem2[3963] = 10'b0010011111;
mem2[3964] = 10'b0010011111;
mem2[3965] = 10'b0010011111;
mem2[3966] = 10'b0010011111;
mem2[3967] = 10'b0010011111;
mem2[3968] = 10'b0010011111;
mem2[3969] = 10'b0010011111;
mem2[3970] = 10'b0010011111;
mem2[3971] = 10'b0010011111;
mem2[3972] = 10'b0010011111;
mem2[3973] = 10'b0010011111;
mem2[3974] = 10'b0010100000;
mem2[3975] = 10'b0010100000;
mem2[3976] = 10'b0010100000;
mem2[3977] = 10'b0010100000;
mem2[3978] = 10'b0010100000;
mem2[3979] = 10'b0010100000;
mem2[3980] = 10'b0010100000;
mem2[3981] = 10'b0010100000;
mem2[3982] = 10'b0010100000;
mem2[3983] = 10'b0010100000;
mem2[3984] = 10'b0010100000;
mem2[3985] = 10'b0010100000;
mem2[3986] = 10'b0010100000;
mem2[3987] = 10'b0010100001;
mem2[3988] = 10'b0010100001;
mem2[3989] = 10'b0010100001;
mem2[3990] = 10'b0010100001;
mem2[3991] = 10'b0010100001;
mem2[3992] = 10'b0010100001;
mem2[3993] = 10'b0010100001;
mem2[3994] = 10'b0010100001;
mem2[3995] = 10'b0010100001;
mem2[3996] = 10'b0010100001;
mem2[3997] = 10'b0010100001;
mem2[3998] = 10'b0010100001;
mem2[3999] = 10'b0010100001;
mem2[4000] = 10'b0010100010;
mem2[4001] = 10'b0010100010;
mem2[4002] = 10'b0010100010;
mem2[4003] = 10'b0010100010;
mem2[4004] = 10'b0010100010;
mem2[4005] = 10'b0010100010;
mem2[4006] = 10'b0010100010;
mem2[4007] = 10'b0010100010;
mem2[4008] = 10'b0010100010;
mem2[4009] = 10'b0010100010;
mem2[4010] = 10'b0010100010;
mem2[4011] = 10'b0010100010;
mem2[4012] = 10'b0010100010;
mem2[4013] = 10'b0010100011;
mem2[4014] = 10'b0010100011;
mem2[4015] = 10'b0010100011;
mem2[4016] = 10'b0010100011;
mem2[4017] = 10'b0010100011;
mem2[4018] = 10'b0010100011;
mem2[4019] = 10'b0010100011;
mem2[4020] = 10'b0010100011;
mem2[4021] = 10'b0010100011;
mem2[4022] = 10'b0010100011;
mem2[4023] = 10'b0010100011;
mem2[4024] = 10'b0010100011;
mem2[4025] = 10'b0010100011;
mem2[4026] = 10'b0010100100;
mem2[4027] = 10'b0010100100;
mem2[4028] = 10'b0010100100;
mem2[4029] = 10'b0010100100;
mem2[4030] = 10'b0010100100;
mem2[4031] = 10'b0010100100;
mem2[4032] = 10'b0010100100;
mem2[4033] = 10'b0010100100;
mem2[4034] = 10'b0010100100;
mem2[4035] = 10'b0010100100;
mem2[4036] = 10'b0010100100;
mem2[4037] = 10'b0010100100;
mem2[4038] = 10'b0010100100;
mem2[4039] = 10'b0010100101;
mem2[4040] = 10'b0010100101;
mem2[4041] = 10'b0010100101;
mem2[4042] = 10'b0010100101;
mem2[4043] = 10'b0010100101;
mem2[4044] = 10'b0010100101;
mem2[4045] = 10'b0010100101;
mem2[4046] = 10'b0010100101;
mem2[4047] = 10'b0010100101;
mem2[4048] = 10'b0010100101;
mem2[4049] = 10'b0010100101;
mem2[4050] = 10'b0010100101;
mem2[4051] = 10'b0010100101;
mem2[4052] = 10'b0010100110;
mem2[4053] = 10'b0010100110;
mem2[4054] = 10'b0010100110;
mem2[4055] = 10'b0010100110;
mem2[4056] = 10'b0010100110;
mem2[4057] = 10'b0010100110;
mem2[4058] = 10'b0010100110;
mem2[4059] = 10'b0010100110;
mem2[4060] = 10'b0010100110;
mem2[4061] = 10'b0010100110;
mem2[4062] = 10'b0010100110;
mem2[4063] = 10'b0010100110;
mem2[4064] = 10'b0010100110;
mem2[4065] = 10'b0010100111;
mem2[4066] = 10'b0010100111;
mem2[4067] = 10'b0010100111;
mem2[4068] = 10'b0010100111;
mem2[4069] = 10'b0010100111;
mem2[4070] = 10'b0010100111;
mem2[4071] = 10'b0010100111;
mem2[4072] = 10'b0010100111;
mem2[4073] = 10'b0010100111;
mem2[4074] = 10'b0010100111;
mem2[4075] = 10'b0010100111;
mem2[4076] = 10'b0010100111;
mem2[4077] = 10'b0010100111;
mem2[4078] = 10'b0010101000;
mem2[4079] = 10'b0010101000;
mem2[4080] = 10'b0010101000;
mem2[4081] = 10'b0010101000;
mem2[4082] = 10'b0010101000;
mem2[4083] = 10'b0010101000;
mem2[4084] = 10'b0010101000;
mem2[4085] = 10'b0010101000;
mem2[4086] = 10'b0010101000;
mem2[4087] = 10'b0010101000;
mem2[4088] = 10'b0010101000;
mem2[4089] = 10'b0010101000;
mem2[4090] = 10'b0010101000;
mem2[4091] = 10'b0010101001;
mem2[4092] = 10'b0010101001;
mem2[4093] = 10'b0010101001;
mem2[4094] = 10'b0010101001;
mem2[4095] = 10'b0010101001;
mem2[4096] = 10'b0010101001;
mem2[4097] = 10'b0010101001;
mem2[4098] = 10'b0010101001;
mem2[4099] = 10'b0010101001;
mem2[4100] = 10'b0010101001;
mem2[4101] = 10'b0010101001;
mem2[4102] = 10'b0010101001;
mem2[4103] = 10'b0010101001;
mem2[4104] = 10'b0010101010;
mem2[4105] = 10'b0010101010;
mem2[4106] = 10'b0010101010;
mem2[4107] = 10'b0010101010;
mem2[4108] = 10'b0010101010;
mem2[4109] = 10'b0010101010;
mem2[4110] = 10'b0010101010;
mem2[4111] = 10'b0010101010;
mem2[4112] = 10'b0010101010;
mem2[4113] = 10'b0010101010;
mem2[4114] = 10'b0010101010;
mem2[4115] = 10'b0010101010;
mem2[4116] = 10'b0010101010;
mem2[4117] = 10'b0010101011;
mem2[4118] = 10'b0010101011;
mem2[4119] = 10'b0010101011;
mem2[4120] = 10'b0010101011;
mem2[4121] = 10'b0010101011;
mem2[4122] = 10'b0010101011;
mem2[4123] = 10'b0010101011;
mem2[4124] = 10'b0010101011;
mem2[4125] = 10'b0010101011;
mem2[4126] = 10'b0010101011;
mem2[4127] = 10'b0010101011;
mem2[4128] = 10'b0010101011;
mem2[4129] = 10'b0010101100;
mem2[4130] = 10'b0010101100;
mem2[4131] = 10'b0010101100;
mem2[4132] = 10'b0010101100;
mem2[4133] = 10'b0010101100;
mem2[4134] = 10'b0010101100;
mem2[4135] = 10'b0010101100;
mem2[4136] = 10'b0010101100;
mem2[4137] = 10'b0010101100;
mem2[4138] = 10'b0010101100;
mem2[4139] = 10'b0010101100;
mem2[4140] = 10'b0010101100;
mem2[4141] = 10'b0010101100;
mem2[4142] = 10'b0010101101;
mem2[4143] = 10'b0010101101;
mem2[4144] = 10'b0010101101;
mem2[4145] = 10'b0010101101;
mem2[4146] = 10'b0010101101;
mem2[4147] = 10'b0010101101;
mem2[4148] = 10'b0010101101;
mem2[4149] = 10'b0010101101;
mem2[4150] = 10'b0010101101;
mem2[4151] = 10'b0010101101;
mem2[4152] = 10'b0010101101;
mem2[4153] = 10'b0010101101;
mem2[4154] = 10'b0010101101;
mem2[4155] = 10'b0010101110;
mem2[4156] = 10'b0010101110;
mem2[4157] = 10'b0010101110;
mem2[4158] = 10'b0010101110;
mem2[4159] = 10'b0010101110;
mem2[4160] = 10'b0010101110;
mem2[4161] = 10'b0010101110;
mem2[4162] = 10'b0010101110;
mem2[4163] = 10'b0010101110;
mem2[4164] = 10'b0010101110;
mem2[4165] = 10'b0010101110;
mem2[4166] = 10'b0010101110;
mem2[4167] = 10'b0010101110;
mem2[4168] = 10'b0010101111;
mem2[4169] = 10'b0010101111;
mem2[4170] = 10'b0010101111;
mem2[4171] = 10'b0010101111;
mem2[4172] = 10'b0010101111;
mem2[4173] = 10'b0010101111;
mem2[4174] = 10'b0010101111;
mem2[4175] = 10'b0010101111;
mem2[4176] = 10'b0010101111;
mem2[4177] = 10'b0010101111;
mem2[4178] = 10'b0010101111;
mem2[4179] = 10'b0010101111;
mem2[4180] = 10'b0010110000;
mem2[4181] = 10'b0010110000;
mem2[4182] = 10'b0010110000;
mem2[4183] = 10'b0010110000;
mem2[4184] = 10'b0010110000;
mem2[4185] = 10'b0010110000;
mem2[4186] = 10'b0010110000;
mem2[4187] = 10'b0010110000;
mem2[4188] = 10'b0010110000;
mem2[4189] = 10'b0010110000;
mem2[4190] = 10'b0010110000;
mem2[4191] = 10'b0010110000;
mem2[4192] = 10'b0010110000;
mem2[4193] = 10'b0010110001;
mem2[4194] = 10'b0010110001;
mem2[4195] = 10'b0010110001;
mem2[4196] = 10'b0010110001;
mem2[4197] = 10'b0010110001;
mem2[4198] = 10'b0010110001;
mem2[4199] = 10'b0010110001;
mem2[4200] = 10'b0010110001;
mem2[4201] = 10'b0010110001;
mem2[4202] = 10'b0010110001;
mem2[4203] = 10'b0010110001;
mem2[4204] = 10'b0010110001;
mem2[4205] = 10'b0010110010;
mem2[4206] = 10'b0010110010;
mem2[4207] = 10'b0010110010;
mem2[4208] = 10'b0010110010;
mem2[4209] = 10'b0010110010;
mem2[4210] = 10'b0010110010;
mem2[4211] = 10'b0010110010;
mem2[4212] = 10'b0010110010;
mem2[4213] = 10'b0010110010;
mem2[4214] = 10'b0010110010;
mem2[4215] = 10'b0010110010;
mem2[4216] = 10'b0010110010;
mem2[4217] = 10'b0010110010;
mem2[4218] = 10'b0010110011;
mem2[4219] = 10'b0010110011;
mem2[4220] = 10'b0010110011;
mem2[4221] = 10'b0010110011;
mem2[4222] = 10'b0010110011;
mem2[4223] = 10'b0010110011;
mem2[4224] = 10'b0010110011;
mem2[4225] = 10'b0010110011;
mem2[4226] = 10'b0010110011;
mem2[4227] = 10'b0010110011;
mem2[4228] = 10'b0010110011;
mem2[4229] = 10'b0010110011;
mem2[4230] = 10'b0010110011;
mem2[4231] = 10'b0010110100;
mem2[4232] = 10'b0010110100;
mem2[4233] = 10'b0010110100;
mem2[4234] = 10'b0010110100;
mem2[4235] = 10'b0010110100;
mem2[4236] = 10'b0010110100;
mem2[4237] = 10'b0010110100;
mem2[4238] = 10'b0010110100;
mem2[4239] = 10'b0010110100;
mem2[4240] = 10'b0010110100;
mem2[4241] = 10'b0010110100;
mem2[4242] = 10'b0010110100;
mem2[4243] = 10'b0010110101;
mem2[4244] = 10'b0010110101;
mem2[4245] = 10'b0010110101;
mem2[4246] = 10'b0010110101;
mem2[4247] = 10'b0010110101;
mem2[4248] = 10'b0010110101;
mem2[4249] = 10'b0010110101;
mem2[4250] = 10'b0010110101;
mem2[4251] = 10'b0010110101;
mem2[4252] = 10'b0010110101;
mem2[4253] = 10'b0010110101;
mem2[4254] = 10'b0010110101;
mem2[4255] = 10'b0010110101;
mem2[4256] = 10'b0010110110;
mem2[4257] = 10'b0010110110;
mem2[4258] = 10'b0010110110;
mem2[4259] = 10'b0010110110;
mem2[4260] = 10'b0010110110;
mem2[4261] = 10'b0010110110;
mem2[4262] = 10'b0010110110;
mem2[4263] = 10'b0010110110;
mem2[4264] = 10'b0010110110;
mem2[4265] = 10'b0010110110;
mem2[4266] = 10'b0010110110;
mem2[4267] = 10'b0010110110;
mem2[4268] = 10'b0010110111;
mem2[4269] = 10'b0010110111;
mem2[4270] = 10'b0010110111;
mem2[4271] = 10'b0010110111;
mem2[4272] = 10'b0010110111;
mem2[4273] = 10'b0010110111;
mem2[4274] = 10'b0010110111;
mem2[4275] = 10'b0010110111;
mem2[4276] = 10'b0010110111;
mem2[4277] = 10'b0010110111;
mem2[4278] = 10'b0010110111;
mem2[4279] = 10'b0010110111;
mem2[4280] = 10'b0010110111;
mem2[4281] = 10'b0010111000;
mem2[4282] = 10'b0010111000;
mem2[4283] = 10'b0010111000;
mem2[4284] = 10'b0010111000;
mem2[4285] = 10'b0010111000;
mem2[4286] = 10'b0010111000;
mem2[4287] = 10'b0010111000;
mem2[4288] = 10'b0010111000;
mem2[4289] = 10'b0010111000;
mem2[4290] = 10'b0010111000;
mem2[4291] = 10'b0010111000;
mem2[4292] = 10'b0010111000;
mem2[4293] = 10'b0010111001;
mem2[4294] = 10'b0010111001;
mem2[4295] = 10'b0010111001;
mem2[4296] = 10'b0010111001;
mem2[4297] = 10'b0010111001;
mem2[4298] = 10'b0010111001;
mem2[4299] = 10'b0010111001;
mem2[4300] = 10'b0010111001;
mem2[4301] = 10'b0010111001;
mem2[4302] = 10'b0010111001;
mem2[4303] = 10'b0010111001;
mem2[4304] = 10'b0010111001;
mem2[4305] = 10'b0010111010;
mem2[4306] = 10'b0010111010;
mem2[4307] = 10'b0010111010;
mem2[4308] = 10'b0010111010;
mem2[4309] = 10'b0010111010;
mem2[4310] = 10'b0010111010;
mem2[4311] = 10'b0010111010;
mem2[4312] = 10'b0010111010;
mem2[4313] = 10'b0010111010;
mem2[4314] = 10'b0010111010;
mem2[4315] = 10'b0010111010;
mem2[4316] = 10'b0010111010;
mem2[4317] = 10'b0010111010;
mem2[4318] = 10'b0010111011;
mem2[4319] = 10'b0010111011;
mem2[4320] = 10'b0010111011;
mem2[4321] = 10'b0010111011;
mem2[4322] = 10'b0010111011;
mem2[4323] = 10'b0010111011;
mem2[4324] = 10'b0010111011;
mem2[4325] = 10'b0010111011;
mem2[4326] = 10'b0010111011;
mem2[4327] = 10'b0010111011;
mem2[4328] = 10'b0010111011;
mem2[4329] = 10'b0010111011;
mem2[4330] = 10'b0010111100;
mem2[4331] = 10'b0010111100;
mem2[4332] = 10'b0010111100;
mem2[4333] = 10'b0010111100;
mem2[4334] = 10'b0010111100;
mem2[4335] = 10'b0010111100;
mem2[4336] = 10'b0010111100;
mem2[4337] = 10'b0010111100;
mem2[4338] = 10'b0010111100;
mem2[4339] = 10'b0010111100;
mem2[4340] = 10'b0010111100;
mem2[4341] = 10'b0010111100;
mem2[4342] = 10'b0010111101;
mem2[4343] = 10'b0010111101;
mem2[4344] = 10'b0010111101;
mem2[4345] = 10'b0010111101;
mem2[4346] = 10'b0010111101;
mem2[4347] = 10'b0010111101;
mem2[4348] = 10'b0010111101;
mem2[4349] = 10'b0010111101;
mem2[4350] = 10'b0010111101;
mem2[4351] = 10'b0010111101;
mem2[4352] = 10'b0010111101;
mem2[4353] = 10'b0010111101;
mem2[4354] = 10'b0010111101;
mem2[4355] = 10'b0010111110;
mem2[4356] = 10'b0010111110;
mem2[4357] = 10'b0010111110;
mem2[4358] = 10'b0010111110;
mem2[4359] = 10'b0010111110;
mem2[4360] = 10'b0010111110;
mem2[4361] = 10'b0010111110;
mem2[4362] = 10'b0010111110;
mem2[4363] = 10'b0010111110;
mem2[4364] = 10'b0010111110;
mem2[4365] = 10'b0010111110;
mem2[4366] = 10'b0010111110;
mem2[4367] = 10'b0010111111;
mem2[4368] = 10'b0010111111;
mem2[4369] = 10'b0010111111;
mem2[4370] = 10'b0010111111;
mem2[4371] = 10'b0010111111;
mem2[4372] = 10'b0010111111;
mem2[4373] = 10'b0010111111;
mem2[4374] = 10'b0010111111;
mem2[4375] = 10'b0010111111;
mem2[4376] = 10'b0010111111;
mem2[4377] = 10'b0010111111;
mem2[4378] = 10'b0010111111;
mem2[4379] = 10'b0011000000;
mem2[4380] = 10'b0011000000;
mem2[4381] = 10'b0011000000;
mem2[4382] = 10'b0011000000;
mem2[4383] = 10'b0011000000;
mem2[4384] = 10'b0011000000;
mem2[4385] = 10'b0011000000;
mem2[4386] = 10'b0011000000;
mem2[4387] = 10'b0011000000;
mem2[4388] = 10'b0011000000;
mem2[4389] = 10'b0011000000;
mem2[4390] = 10'b0011000000;
mem2[4391] = 10'b0011000001;
mem2[4392] = 10'b0011000001;
mem2[4393] = 10'b0011000001;
mem2[4394] = 10'b0011000001;
mem2[4395] = 10'b0011000001;
mem2[4396] = 10'b0011000001;
mem2[4397] = 10'b0011000001;
mem2[4398] = 10'b0011000001;
mem2[4399] = 10'b0011000001;
mem2[4400] = 10'b0011000001;
mem2[4401] = 10'b0011000001;
mem2[4402] = 10'b0011000001;
mem2[4403] = 10'b0011000001;
mem2[4404] = 10'b0011000010;
mem2[4405] = 10'b0011000010;
mem2[4406] = 10'b0011000010;
mem2[4407] = 10'b0011000010;
mem2[4408] = 10'b0011000010;
mem2[4409] = 10'b0011000010;
mem2[4410] = 10'b0011000010;
mem2[4411] = 10'b0011000010;
mem2[4412] = 10'b0011000010;
mem2[4413] = 10'b0011000010;
mem2[4414] = 10'b0011000010;
mem2[4415] = 10'b0011000010;
mem2[4416] = 10'b0011000011;
mem2[4417] = 10'b0011000011;
mem2[4418] = 10'b0011000011;
mem2[4419] = 10'b0011000011;
mem2[4420] = 10'b0011000011;
mem2[4421] = 10'b0011000011;
mem2[4422] = 10'b0011000011;
mem2[4423] = 10'b0011000011;
mem2[4424] = 10'b0011000011;
mem2[4425] = 10'b0011000011;
mem2[4426] = 10'b0011000011;
mem2[4427] = 10'b0011000011;
mem2[4428] = 10'b0011000100;
mem2[4429] = 10'b0011000100;
mem2[4430] = 10'b0011000100;
mem2[4431] = 10'b0011000100;
mem2[4432] = 10'b0011000100;
mem2[4433] = 10'b0011000100;
mem2[4434] = 10'b0011000100;
mem2[4435] = 10'b0011000100;
mem2[4436] = 10'b0011000100;
mem2[4437] = 10'b0011000100;
mem2[4438] = 10'b0011000100;
mem2[4439] = 10'b0011000100;
mem2[4440] = 10'b0011000101;
mem2[4441] = 10'b0011000101;
mem2[4442] = 10'b0011000101;
mem2[4443] = 10'b0011000101;
mem2[4444] = 10'b0011000101;
mem2[4445] = 10'b0011000101;
mem2[4446] = 10'b0011000101;
mem2[4447] = 10'b0011000101;
mem2[4448] = 10'b0011000101;
mem2[4449] = 10'b0011000101;
mem2[4450] = 10'b0011000101;
mem2[4451] = 10'b0011000101;
mem2[4452] = 10'b0011000110;
mem2[4453] = 10'b0011000110;
mem2[4454] = 10'b0011000110;
mem2[4455] = 10'b0011000110;
mem2[4456] = 10'b0011000110;
mem2[4457] = 10'b0011000110;
mem2[4458] = 10'b0011000110;
mem2[4459] = 10'b0011000110;
mem2[4460] = 10'b0011000110;
mem2[4461] = 10'b0011000110;
mem2[4462] = 10'b0011000110;
mem2[4463] = 10'b0011000110;
mem2[4464] = 10'b0011000111;
mem2[4465] = 10'b0011000111;
mem2[4466] = 10'b0011000111;
mem2[4467] = 10'b0011000111;
mem2[4468] = 10'b0011000111;
mem2[4469] = 10'b0011000111;
mem2[4470] = 10'b0011000111;
mem2[4471] = 10'b0011000111;
mem2[4472] = 10'b0011000111;
mem2[4473] = 10'b0011000111;
mem2[4474] = 10'b0011000111;
mem2[4475] = 10'b0011000111;
mem2[4476] = 10'b0011001000;
mem2[4477] = 10'b0011001000;
mem2[4478] = 10'b0011001000;
mem2[4479] = 10'b0011001000;
mem2[4480] = 10'b0011001000;
mem2[4481] = 10'b0011001000;
mem2[4482] = 10'b0011001000;
mem2[4483] = 10'b0011001000;
mem2[4484] = 10'b0011001000;
mem2[4485] = 10'b0011001000;
mem2[4486] = 10'b0011001000;
mem2[4487] = 10'b0011001000;
mem2[4488] = 10'b0011001001;
mem2[4489] = 10'b0011001001;
mem2[4490] = 10'b0011001001;
mem2[4491] = 10'b0011001001;
mem2[4492] = 10'b0011001001;
mem2[4493] = 10'b0011001001;
mem2[4494] = 10'b0011001001;
mem2[4495] = 10'b0011001001;
mem2[4496] = 10'b0011001001;
mem2[4497] = 10'b0011001001;
mem2[4498] = 10'b0011001001;
mem2[4499] = 10'b0011001001;
mem2[4500] = 10'b0011001010;
mem2[4501] = 10'b0011001010;
mem2[4502] = 10'b0011001010;
mem2[4503] = 10'b0011001010;
mem2[4504] = 10'b0011001010;
mem2[4505] = 10'b0011001010;
mem2[4506] = 10'b0011001010;
mem2[4507] = 10'b0011001010;
mem2[4508] = 10'b0011001010;
mem2[4509] = 10'b0011001010;
mem2[4510] = 10'b0011001010;
mem2[4511] = 10'b0011001010;
mem2[4512] = 10'b0011001011;
mem2[4513] = 10'b0011001011;
mem2[4514] = 10'b0011001011;
mem2[4515] = 10'b0011001011;
mem2[4516] = 10'b0011001011;
mem2[4517] = 10'b0011001011;
mem2[4518] = 10'b0011001011;
mem2[4519] = 10'b0011001011;
mem2[4520] = 10'b0011001011;
mem2[4521] = 10'b0011001011;
mem2[4522] = 10'b0011001011;
mem2[4523] = 10'b0011001011;
mem2[4524] = 10'b0011001100;
mem2[4525] = 10'b0011001100;
mem2[4526] = 10'b0011001100;
mem2[4527] = 10'b0011001100;
mem2[4528] = 10'b0011001100;
mem2[4529] = 10'b0011001100;
mem2[4530] = 10'b0011001100;
mem2[4531] = 10'b0011001100;
mem2[4532] = 10'b0011001100;
mem2[4533] = 10'b0011001100;
mem2[4534] = 10'b0011001100;
mem2[4535] = 10'b0011001100;
mem2[4536] = 10'b0011001101;
mem2[4537] = 10'b0011001101;
mem2[4538] = 10'b0011001101;
mem2[4539] = 10'b0011001101;
mem2[4540] = 10'b0011001101;
mem2[4541] = 10'b0011001101;
mem2[4542] = 10'b0011001101;
mem2[4543] = 10'b0011001101;
mem2[4544] = 10'b0011001101;
mem2[4545] = 10'b0011001101;
mem2[4546] = 10'b0011001101;
mem2[4547] = 10'b0011001101;
mem2[4548] = 10'b0011001110;
mem2[4549] = 10'b0011001110;
mem2[4550] = 10'b0011001110;
mem2[4551] = 10'b0011001110;
mem2[4552] = 10'b0011001110;
mem2[4553] = 10'b0011001110;
mem2[4554] = 10'b0011001110;
mem2[4555] = 10'b0011001110;
mem2[4556] = 10'b0011001110;
mem2[4557] = 10'b0011001110;
mem2[4558] = 10'b0011001110;
mem2[4559] = 10'b0011001110;
mem2[4560] = 10'b0011001111;
mem2[4561] = 10'b0011001111;
mem2[4562] = 10'b0011001111;
mem2[4563] = 10'b0011001111;
mem2[4564] = 10'b0011001111;
mem2[4565] = 10'b0011001111;
mem2[4566] = 10'b0011001111;
mem2[4567] = 10'b0011001111;
mem2[4568] = 10'b0011001111;
mem2[4569] = 10'b0011001111;
mem2[4570] = 10'b0011001111;
mem2[4571] = 10'b0011001111;
mem2[4572] = 10'b0011010000;
mem2[4573] = 10'b0011010000;
mem2[4574] = 10'b0011010000;
mem2[4575] = 10'b0011010000;
mem2[4576] = 10'b0011010000;
mem2[4577] = 10'b0011010000;
mem2[4578] = 10'b0011010000;
mem2[4579] = 10'b0011010000;
mem2[4580] = 10'b0011010000;
mem2[4581] = 10'b0011010000;
mem2[4582] = 10'b0011010000;
mem2[4583] = 10'b0011010000;
mem2[4584] = 10'b0011010001;
mem2[4585] = 10'b0011010001;
mem2[4586] = 10'b0011010001;
mem2[4587] = 10'b0011010001;
mem2[4588] = 10'b0011010001;
mem2[4589] = 10'b0011010001;
mem2[4590] = 10'b0011010001;
mem2[4591] = 10'b0011010001;
mem2[4592] = 10'b0011010001;
mem2[4593] = 10'b0011010001;
mem2[4594] = 10'b0011010001;
mem2[4595] = 10'b0011010001;
mem2[4596] = 10'b0011010010;
mem2[4597] = 10'b0011010010;
mem2[4598] = 10'b0011010010;
mem2[4599] = 10'b0011010010;
mem2[4600] = 10'b0011010010;
mem2[4601] = 10'b0011010010;
mem2[4602] = 10'b0011010010;
mem2[4603] = 10'b0011010010;
mem2[4604] = 10'b0011010010;
mem2[4605] = 10'b0011010010;
mem2[4606] = 10'b0011010010;
mem2[4607] = 10'b0011010011;
mem2[4608] = 10'b0011010011;
mem2[4609] = 10'b0011010011;
mem2[4610] = 10'b0011010011;
mem2[4611] = 10'b0011010011;
mem2[4612] = 10'b0011010011;
mem2[4613] = 10'b0011010011;
mem2[4614] = 10'b0011010011;
mem2[4615] = 10'b0011010011;
mem2[4616] = 10'b0011010011;
mem2[4617] = 10'b0011010011;
mem2[4618] = 10'b0011010011;
mem2[4619] = 10'b0011010100;
mem2[4620] = 10'b0011010100;
mem2[4621] = 10'b0011010100;
mem2[4622] = 10'b0011010100;
mem2[4623] = 10'b0011010100;
mem2[4624] = 10'b0011010100;
mem2[4625] = 10'b0011010100;
mem2[4626] = 10'b0011010100;
mem2[4627] = 10'b0011010100;
mem2[4628] = 10'b0011010100;
mem2[4629] = 10'b0011010100;
mem2[4630] = 10'b0011010100;
mem2[4631] = 10'b0011010101;
mem2[4632] = 10'b0011010101;
mem2[4633] = 10'b0011010101;
mem2[4634] = 10'b0011010101;
mem2[4635] = 10'b0011010101;
mem2[4636] = 10'b0011010101;
mem2[4637] = 10'b0011010101;
mem2[4638] = 10'b0011010101;
mem2[4639] = 10'b0011010101;
mem2[4640] = 10'b0011010101;
mem2[4641] = 10'b0011010101;
mem2[4642] = 10'b0011010101;
mem2[4643] = 10'b0011010110;
mem2[4644] = 10'b0011010110;
mem2[4645] = 10'b0011010110;
mem2[4646] = 10'b0011010110;
mem2[4647] = 10'b0011010110;
mem2[4648] = 10'b0011010110;
mem2[4649] = 10'b0011010110;
mem2[4650] = 10'b0011010110;
mem2[4651] = 10'b0011010110;
mem2[4652] = 10'b0011010110;
mem2[4653] = 10'b0011010110;
mem2[4654] = 10'b0011010110;
mem2[4655] = 10'b0011010111;
mem2[4656] = 10'b0011010111;
mem2[4657] = 10'b0011010111;
mem2[4658] = 10'b0011010111;
mem2[4659] = 10'b0011010111;
mem2[4660] = 10'b0011010111;
mem2[4661] = 10'b0011010111;
mem2[4662] = 10'b0011010111;
mem2[4663] = 10'b0011010111;
mem2[4664] = 10'b0011010111;
mem2[4665] = 10'b0011010111;
mem2[4666] = 10'b0011011000;
mem2[4667] = 10'b0011011000;
mem2[4668] = 10'b0011011000;
mem2[4669] = 10'b0011011000;
mem2[4670] = 10'b0011011000;
mem2[4671] = 10'b0011011000;
mem2[4672] = 10'b0011011000;
mem2[4673] = 10'b0011011000;
mem2[4674] = 10'b0011011000;
mem2[4675] = 10'b0011011000;
mem2[4676] = 10'b0011011000;
mem2[4677] = 10'b0011011000;
mem2[4678] = 10'b0011011001;
mem2[4679] = 10'b0011011001;
mem2[4680] = 10'b0011011001;
mem2[4681] = 10'b0011011001;
mem2[4682] = 10'b0011011001;
mem2[4683] = 10'b0011011001;
mem2[4684] = 10'b0011011001;
mem2[4685] = 10'b0011011001;
mem2[4686] = 10'b0011011001;
mem2[4687] = 10'b0011011001;
mem2[4688] = 10'b0011011001;
mem2[4689] = 10'b0011011001;
mem2[4690] = 10'b0011011010;
mem2[4691] = 10'b0011011010;
mem2[4692] = 10'b0011011010;
mem2[4693] = 10'b0011011010;
mem2[4694] = 10'b0011011010;
mem2[4695] = 10'b0011011010;
mem2[4696] = 10'b0011011010;
mem2[4697] = 10'b0011011010;
mem2[4698] = 10'b0011011010;
mem2[4699] = 10'b0011011010;
mem2[4700] = 10'b0011011010;
mem2[4701] = 10'b0011011011;
mem2[4702] = 10'b0011011011;
mem2[4703] = 10'b0011011011;
mem2[4704] = 10'b0011011011;
mem2[4705] = 10'b0011011011;
mem2[4706] = 10'b0011011011;
mem2[4707] = 10'b0011011011;
mem2[4708] = 10'b0011011011;
mem2[4709] = 10'b0011011011;
mem2[4710] = 10'b0011011011;
mem2[4711] = 10'b0011011011;
mem2[4712] = 10'b0011011011;
mem2[4713] = 10'b0011011100;
mem2[4714] = 10'b0011011100;
mem2[4715] = 10'b0011011100;
mem2[4716] = 10'b0011011100;
mem2[4717] = 10'b0011011100;
mem2[4718] = 10'b0011011100;
mem2[4719] = 10'b0011011100;
mem2[4720] = 10'b0011011100;
mem2[4721] = 10'b0011011100;
mem2[4722] = 10'b0011011100;
mem2[4723] = 10'b0011011100;
mem2[4724] = 10'b0011011101;
mem2[4725] = 10'b0011011101;
mem2[4726] = 10'b0011011101;
mem2[4727] = 10'b0011011101;
mem2[4728] = 10'b0011011101;
mem2[4729] = 10'b0011011101;
mem2[4730] = 10'b0011011101;
mem2[4731] = 10'b0011011101;
mem2[4732] = 10'b0011011101;
mem2[4733] = 10'b0011011101;
mem2[4734] = 10'b0011011101;
mem2[4735] = 10'b0011011101;
mem2[4736] = 10'b0011011110;
mem2[4737] = 10'b0011011110;
mem2[4738] = 10'b0011011110;
mem2[4739] = 10'b0011011110;
mem2[4740] = 10'b0011011110;
mem2[4741] = 10'b0011011110;
mem2[4742] = 10'b0011011110;
mem2[4743] = 10'b0011011110;
mem2[4744] = 10'b0011011110;
mem2[4745] = 10'b0011011110;
mem2[4746] = 10'b0011011110;
mem2[4747] = 10'b0011011110;
mem2[4748] = 10'b0011011111;
mem2[4749] = 10'b0011011111;
mem2[4750] = 10'b0011011111;
mem2[4751] = 10'b0011011111;
mem2[4752] = 10'b0011011111;
mem2[4753] = 10'b0011011111;
mem2[4754] = 10'b0011011111;
mem2[4755] = 10'b0011011111;
mem2[4756] = 10'b0011011111;
mem2[4757] = 10'b0011011111;
mem2[4758] = 10'b0011011111;
mem2[4759] = 10'b0011100000;
mem2[4760] = 10'b0011100000;
mem2[4761] = 10'b0011100000;
mem2[4762] = 10'b0011100000;
mem2[4763] = 10'b0011100000;
mem2[4764] = 10'b0011100000;
mem2[4765] = 10'b0011100000;
mem2[4766] = 10'b0011100000;
mem2[4767] = 10'b0011100000;
mem2[4768] = 10'b0011100000;
mem2[4769] = 10'b0011100000;
mem2[4770] = 10'b0011100000;
mem2[4771] = 10'b0011100001;
mem2[4772] = 10'b0011100001;
mem2[4773] = 10'b0011100001;
mem2[4774] = 10'b0011100001;
mem2[4775] = 10'b0011100001;
mem2[4776] = 10'b0011100001;
mem2[4777] = 10'b0011100001;
mem2[4778] = 10'b0011100001;
mem2[4779] = 10'b0011100001;
mem2[4780] = 10'b0011100001;
mem2[4781] = 10'b0011100001;
mem2[4782] = 10'b0011100010;
mem2[4783] = 10'b0011100010;
mem2[4784] = 10'b0011100010;
mem2[4785] = 10'b0011100010;
mem2[4786] = 10'b0011100010;
mem2[4787] = 10'b0011100010;
mem2[4788] = 10'b0011100010;
mem2[4789] = 10'b0011100010;
mem2[4790] = 10'b0011100010;
mem2[4791] = 10'b0011100010;
mem2[4792] = 10'b0011100010;
mem2[4793] = 10'b0011100010;
mem2[4794] = 10'b0011100011;
mem2[4795] = 10'b0011100011;
mem2[4796] = 10'b0011100011;
mem2[4797] = 10'b0011100011;
mem2[4798] = 10'b0011100011;
mem2[4799] = 10'b0011100011;
mem2[4800] = 10'b0011100011;
mem2[4801] = 10'b0011100011;
mem2[4802] = 10'b0011100011;
mem2[4803] = 10'b0011100011;
mem2[4804] = 10'b0011100011;
mem2[4805] = 10'b0011100100;
mem2[4806] = 10'b0011100100;
mem2[4807] = 10'b0011100100;
mem2[4808] = 10'b0011100100;
mem2[4809] = 10'b0011100100;
mem2[4810] = 10'b0011100100;
mem2[4811] = 10'b0011100100;
mem2[4812] = 10'b0011100100;
mem2[4813] = 10'b0011100100;
mem2[4814] = 10'b0011100100;
mem2[4815] = 10'b0011100100;
mem2[4816] = 10'b0011100100;
mem2[4817] = 10'b0011100101;
mem2[4818] = 10'b0011100101;
mem2[4819] = 10'b0011100101;
mem2[4820] = 10'b0011100101;
mem2[4821] = 10'b0011100101;
mem2[4822] = 10'b0011100101;
mem2[4823] = 10'b0011100101;
mem2[4824] = 10'b0011100101;
mem2[4825] = 10'b0011100101;
mem2[4826] = 10'b0011100101;
mem2[4827] = 10'b0011100101;
mem2[4828] = 10'b0011100110;
mem2[4829] = 10'b0011100110;
mem2[4830] = 10'b0011100110;
mem2[4831] = 10'b0011100110;
mem2[4832] = 10'b0011100110;
mem2[4833] = 10'b0011100110;
mem2[4834] = 10'b0011100110;
mem2[4835] = 10'b0011100110;
mem2[4836] = 10'b0011100110;
mem2[4837] = 10'b0011100110;
mem2[4838] = 10'b0011100110;
mem2[4839] = 10'b0011100110;
mem2[4840] = 10'b0011100111;
mem2[4841] = 10'b0011100111;
mem2[4842] = 10'b0011100111;
mem2[4843] = 10'b0011100111;
mem2[4844] = 10'b0011100111;
mem2[4845] = 10'b0011100111;
mem2[4846] = 10'b0011100111;
mem2[4847] = 10'b0011100111;
mem2[4848] = 10'b0011100111;
mem2[4849] = 10'b0011100111;
mem2[4850] = 10'b0011100111;
mem2[4851] = 10'b0011101000;
mem2[4852] = 10'b0011101000;
mem2[4853] = 10'b0011101000;
mem2[4854] = 10'b0011101000;
mem2[4855] = 10'b0011101000;
mem2[4856] = 10'b0011101000;
mem2[4857] = 10'b0011101000;
mem2[4858] = 10'b0011101000;
mem2[4859] = 10'b0011101000;
mem2[4860] = 10'b0011101000;
mem2[4861] = 10'b0011101000;
mem2[4862] = 10'b0011101001;
mem2[4863] = 10'b0011101001;
mem2[4864] = 10'b0011101001;
mem2[4865] = 10'b0011101001;
mem2[4866] = 10'b0011101001;
mem2[4867] = 10'b0011101001;
mem2[4868] = 10'b0011101001;
mem2[4869] = 10'b0011101001;
mem2[4870] = 10'b0011101001;
mem2[4871] = 10'b0011101001;
mem2[4872] = 10'b0011101001;
mem2[4873] = 10'b0011101001;
mem2[4874] = 10'b0011101010;
mem2[4875] = 10'b0011101010;
mem2[4876] = 10'b0011101010;
mem2[4877] = 10'b0011101010;
mem2[4878] = 10'b0011101010;
mem2[4879] = 10'b0011101010;
mem2[4880] = 10'b0011101010;
mem2[4881] = 10'b0011101010;
mem2[4882] = 10'b0011101010;
mem2[4883] = 10'b0011101010;
mem2[4884] = 10'b0011101010;
mem2[4885] = 10'b0011101011;
mem2[4886] = 10'b0011101011;
mem2[4887] = 10'b0011101011;
mem2[4888] = 10'b0011101011;
mem2[4889] = 10'b0011101011;
mem2[4890] = 10'b0011101011;
mem2[4891] = 10'b0011101011;
mem2[4892] = 10'b0011101011;
mem2[4893] = 10'b0011101011;
mem2[4894] = 10'b0011101011;
mem2[4895] = 10'b0011101011;
mem2[4896] = 10'b0011101011;
mem2[4897] = 10'b0011101100;
mem2[4898] = 10'b0011101100;
mem2[4899] = 10'b0011101100;
mem2[4900] = 10'b0011101100;
mem2[4901] = 10'b0011101100;
mem2[4902] = 10'b0011101100;
mem2[4903] = 10'b0011101100;
mem2[4904] = 10'b0011101100;
mem2[4905] = 10'b0011101100;
mem2[4906] = 10'b0011101100;
mem2[4907] = 10'b0011101100;
mem2[4908] = 10'b0011101101;
mem2[4909] = 10'b0011101101;
mem2[4910] = 10'b0011101101;
mem2[4911] = 10'b0011101101;
mem2[4912] = 10'b0011101101;
mem2[4913] = 10'b0011101101;
mem2[4914] = 10'b0011101101;
mem2[4915] = 10'b0011101101;
mem2[4916] = 10'b0011101101;
mem2[4917] = 10'b0011101101;
mem2[4918] = 10'b0011101101;
mem2[4919] = 10'b0011101110;
mem2[4920] = 10'b0011101110;
mem2[4921] = 10'b0011101110;
mem2[4922] = 10'b0011101110;
mem2[4923] = 10'b0011101110;
mem2[4924] = 10'b0011101110;
mem2[4925] = 10'b0011101110;
mem2[4926] = 10'b0011101110;
mem2[4927] = 10'b0011101110;
mem2[4928] = 10'b0011101110;
mem2[4929] = 10'b0011101110;
mem2[4930] = 10'b0011101111;
mem2[4931] = 10'b0011101111;
mem2[4932] = 10'b0011101111;
mem2[4933] = 10'b0011101111;
mem2[4934] = 10'b0011101111;
mem2[4935] = 10'b0011101111;
mem2[4936] = 10'b0011101111;
mem2[4937] = 10'b0011101111;
mem2[4938] = 10'b0011101111;
mem2[4939] = 10'b0011101111;
mem2[4940] = 10'b0011101111;
mem2[4941] = 10'b0011101111;
mem2[4942] = 10'b0011110000;
mem2[4943] = 10'b0011110000;
mem2[4944] = 10'b0011110000;
mem2[4945] = 10'b0011110000;
mem2[4946] = 10'b0011110000;
mem2[4947] = 10'b0011110000;
mem2[4948] = 10'b0011110000;
mem2[4949] = 10'b0011110000;
mem2[4950] = 10'b0011110000;
mem2[4951] = 10'b0011110000;
mem2[4952] = 10'b0011110000;
mem2[4953] = 10'b0011110001;
mem2[4954] = 10'b0011110001;
mem2[4955] = 10'b0011110001;
mem2[4956] = 10'b0011110001;
mem2[4957] = 10'b0011110001;
mem2[4958] = 10'b0011110001;
mem2[4959] = 10'b0011110001;
mem2[4960] = 10'b0011110001;
mem2[4961] = 10'b0011110001;
mem2[4962] = 10'b0011110001;
mem2[4963] = 10'b0011110001;
mem2[4964] = 10'b0011110010;
mem2[4965] = 10'b0011110010;
mem2[4966] = 10'b0011110010;
mem2[4967] = 10'b0011110010;
mem2[4968] = 10'b0011110010;
mem2[4969] = 10'b0011110010;
mem2[4970] = 10'b0011110010;
mem2[4971] = 10'b0011110010;
mem2[4972] = 10'b0011110010;
mem2[4973] = 10'b0011110010;
mem2[4974] = 10'b0011110010;
mem2[4975] = 10'b0011110011;
mem2[4976] = 10'b0011110011;
mem2[4977] = 10'b0011110011;
mem2[4978] = 10'b0011110011;
mem2[4979] = 10'b0011110011;
mem2[4980] = 10'b0011110011;
mem2[4981] = 10'b0011110011;
mem2[4982] = 10'b0011110011;
mem2[4983] = 10'b0011110011;
mem2[4984] = 10'b0011110011;
mem2[4985] = 10'b0011110011;
mem2[4986] = 10'b0011110011;
mem2[4987] = 10'b0011110100;
mem2[4988] = 10'b0011110100;
mem2[4989] = 10'b0011110100;
mem2[4990] = 10'b0011110100;
mem2[4991] = 10'b0011110100;
mem2[4992] = 10'b0011110100;
mem2[4993] = 10'b0011110100;
mem2[4994] = 10'b0011110100;
mem2[4995] = 10'b0011110100;
mem2[4996] = 10'b0011110100;
mem2[4997] = 10'b0011110100;
mem2[4998] = 10'b0011110101;
mem2[4999] = 10'b0011110101;
mem2[5000] = 10'b0011110101;
mem2[5001] = 10'b0011110101;
mem2[5002] = 10'b0011110101;
mem2[5003] = 10'b0011110101;
mem2[5004] = 10'b0011110101;
mem2[5005] = 10'b0011110101;
mem2[5006] = 10'b0011110101;
mem2[5007] = 10'b0011110101;
mem2[5008] = 10'b0011110101;
mem2[5009] = 10'b0011110110;
mem2[5010] = 10'b0011110110;
mem2[5011] = 10'b0011110110;
mem2[5012] = 10'b0011110110;
mem2[5013] = 10'b0011110110;
mem2[5014] = 10'b0011110110;
mem2[5015] = 10'b0011110110;
mem2[5016] = 10'b0011110110;
mem2[5017] = 10'b0011110110;
mem2[5018] = 10'b0011110110;
mem2[5019] = 10'b0011110110;
mem2[5020] = 10'b0011110111;
mem2[5021] = 10'b0011110111;
mem2[5022] = 10'b0011110111;
mem2[5023] = 10'b0011110111;
mem2[5024] = 10'b0011110111;
mem2[5025] = 10'b0011110111;
mem2[5026] = 10'b0011110111;
mem2[5027] = 10'b0011110111;
mem2[5028] = 10'b0011110111;
mem2[5029] = 10'b0011110111;
mem2[5030] = 10'b0011110111;
mem2[5031] = 10'b0011111000;
mem2[5032] = 10'b0011111000;
mem2[5033] = 10'b0011111000;
mem2[5034] = 10'b0011111000;
mem2[5035] = 10'b0011111000;
mem2[5036] = 10'b0011111000;
mem2[5037] = 10'b0011111000;
mem2[5038] = 10'b0011111000;
mem2[5039] = 10'b0011111000;
mem2[5040] = 10'b0011111000;
mem2[5041] = 10'b0011111000;
mem2[5042] = 10'b0011111000;
mem2[5043] = 10'b0011111001;
mem2[5044] = 10'b0011111001;
mem2[5045] = 10'b0011111001;
mem2[5046] = 10'b0011111001;
mem2[5047] = 10'b0011111001;
mem2[5048] = 10'b0011111001;
mem2[5049] = 10'b0011111001;
mem2[5050] = 10'b0011111001;
mem2[5051] = 10'b0011111001;
mem2[5052] = 10'b0011111001;
mem2[5053] = 10'b0011111001;
mem2[5054] = 10'b0011111010;
mem2[5055] = 10'b0011111010;
mem2[5056] = 10'b0011111010;
mem2[5057] = 10'b0011111010;
mem2[5058] = 10'b0011111010;
mem2[5059] = 10'b0011111010;
mem2[5060] = 10'b0011111010;
mem2[5061] = 10'b0011111010;
mem2[5062] = 10'b0011111010;
mem2[5063] = 10'b0011111010;
mem2[5064] = 10'b0011111010;
mem2[5065] = 10'b0011111011;
mem2[5066] = 10'b0011111011;
mem2[5067] = 10'b0011111011;
mem2[5068] = 10'b0011111011;
mem2[5069] = 10'b0011111011;
mem2[5070] = 10'b0011111011;
mem2[5071] = 10'b0011111011;
mem2[5072] = 10'b0011111011;
mem2[5073] = 10'b0011111011;
mem2[5074] = 10'b0011111011;
mem2[5075] = 10'b0011111011;
mem2[5076] = 10'b0011111100;
mem2[5077] = 10'b0011111100;
mem2[5078] = 10'b0011111100;
mem2[5079] = 10'b0011111100;
mem2[5080] = 10'b0011111100;
mem2[5081] = 10'b0011111100;
mem2[5082] = 10'b0011111100;
mem2[5083] = 10'b0011111100;
mem2[5084] = 10'b0011111100;
mem2[5085] = 10'b0011111100;
mem2[5086] = 10'b0011111100;
mem2[5087] = 10'b0011111101;
mem2[5088] = 10'b0011111101;
mem2[5089] = 10'b0011111101;
mem2[5090] = 10'b0011111101;
mem2[5091] = 10'b0011111101;
mem2[5092] = 10'b0011111101;
mem2[5093] = 10'b0011111101;
mem2[5094] = 10'b0011111101;
mem2[5095] = 10'b0011111101;
mem2[5096] = 10'b0011111101;
mem2[5097] = 10'b0011111101;
mem2[5098] = 10'b0011111110;
mem2[5099] = 10'b0011111110;
mem2[5100] = 10'b0011111110;
mem2[5101] = 10'b0011111110;
mem2[5102] = 10'b0011111110;
mem2[5103] = 10'b0011111110;
mem2[5104] = 10'b0011111110;
mem2[5105] = 10'b0011111110;
mem2[5106] = 10'b0011111110;
mem2[5107] = 10'b0011111110;
mem2[5108] = 10'b0011111110;
mem2[5109] = 10'b0011111111;
mem2[5110] = 10'b0011111111;
mem2[5111] = 10'b0011111111;
mem2[5112] = 10'b0011111111;
mem2[5113] = 10'b0011111111;
mem2[5114] = 10'b0011111111;
mem2[5115] = 10'b0011111111;
mem2[5116] = 10'b0011111111;
mem2[5117] = 10'b0011111111;
mem2[5118] = 10'b0011111111;
mem2[5119] = 10'b0011111111;
mem2[5120] = 10'b0100000000;
mem2[5121] = 10'b0100000000;
mem2[5122] = 10'b0100000000;
mem2[5123] = 10'b0100000000;
mem2[5124] = 10'b0100000000;
mem2[5125] = 10'b0100000000;
mem2[5126] = 10'b0100000000;
mem2[5127] = 10'b0100000000;
mem2[5128] = 10'b0100000000;
mem2[5129] = 10'b0100000000;
mem2[5130] = 10'b0100000000;
mem2[5131] = 10'b0100000001;
mem2[5132] = 10'b0100000001;
mem2[5133] = 10'b0100000001;
mem2[5134] = 10'b0100000001;
mem2[5135] = 10'b0100000001;
mem2[5136] = 10'b0100000001;
mem2[5137] = 10'b0100000001;
mem2[5138] = 10'b0100000001;
mem2[5139] = 10'b0100000001;
mem2[5140] = 10'b0100000001;
mem2[5141] = 10'b0100000001;
mem2[5142] = 10'b0100000010;
mem2[5143] = 10'b0100000010;
mem2[5144] = 10'b0100000010;
mem2[5145] = 10'b0100000010;
mem2[5146] = 10'b0100000010;
mem2[5147] = 10'b0100000010;
mem2[5148] = 10'b0100000010;
mem2[5149] = 10'b0100000010;
mem2[5150] = 10'b0100000010;
mem2[5151] = 10'b0100000010;
mem2[5152] = 10'b0100000010;
mem2[5153] = 10'b0100000011;
mem2[5154] = 10'b0100000011;
mem2[5155] = 10'b0100000011;
mem2[5156] = 10'b0100000011;
mem2[5157] = 10'b0100000011;
mem2[5158] = 10'b0100000011;
mem2[5159] = 10'b0100000011;
mem2[5160] = 10'b0100000011;
mem2[5161] = 10'b0100000011;
mem2[5162] = 10'b0100000011;
mem2[5163] = 10'b0100000011;
mem2[5164] = 10'b0100000100;
mem2[5165] = 10'b0100000100;
mem2[5166] = 10'b0100000100;
mem2[5167] = 10'b0100000100;
mem2[5168] = 10'b0100000100;
mem2[5169] = 10'b0100000100;
mem2[5170] = 10'b0100000100;
mem2[5171] = 10'b0100000100;
mem2[5172] = 10'b0100000100;
mem2[5173] = 10'b0100000100;
mem2[5174] = 10'b0100000100;
mem2[5175] = 10'b0100000101;
mem2[5176] = 10'b0100000101;
mem2[5177] = 10'b0100000101;
mem2[5178] = 10'b0100000101;
mem2[5179] = 10'b0100000101;
mem2[5180] = 10'b0100000101;
mem2[5181] = 10'b0100000101;
mem2[5182] = 10'b0100000101;
mem2[5183] = 10'b0100000101;
mem2[5184] = 10'b0100000101;
mem2[5185] = 10'b0100000101;
mem2[5186] = 10'b0100000110;
mem2[5187] = 10'b0100000110;
mem2[5188] = 10'b0100000110;
mem2[5189] = 10'b0100000110;
mem2[5190] = 10'b0100000110;
mem2[5191] = 10'b0100000110;
mem2[5192] = 10'b0100000110;
mem2[5193] = 10'b0100000110;
mem2[5194] = 10'b0100000110;
mem2[5195] = 10'b0100000110;
mem2[5196] = 10'b0100000110;
mem2[5197] = 10'b0100000111;
mem2[5198] = 10'b0100000111;
mem2[5199] = 10'b0100000111;
mem2[5200] = 10'b0100000111;
mem2[5201] = 10'b0100000111;
mem2[5202] = 10'b0100000111;
mem2[5203] = 10'b0100000111;
mem2[5204] = 10'b0100000111;
mem2[5205] = 10'b0100000111;
mem2[5206] = 10'b0100000111;
mem2[5207] = 10'b0100000111;
mem2[5208] = 10'b0100001000;
mem2[5209] = 10'b0100001000;
mem2[5210] = 10'b0100001000;
mem2[5211] = 10'b0100001000;
mem2[5212] = 10'b0100001000;
mem2[5213] = 10'b0100001000;
mem2[5214] = 10'b0100001000;
mem2[5215] = 10'b0100001000;
mem2[5216] = 10'b0100001000;
mem2[5217] = 10'b0100001000;
mem2[5218] = 10'b0100001000;
mem2[5219] = 10'b0100001001;
mem2[5220] = 10'b0100001001;
mem2[5221] = 10'b0100001001;
mem2[5222] = 10'b0100001001;
mem2[5223] = 10'b0100001001;
mem2[5224] = 10'b0100001001;
mem2[5225] = 10'b0100001001;
mem2[5226] = 10'b0100001001;
mem2[5227] = 10'b0100001001;
mem2[5228] = 10'b0100001001;
mem2[5229] = 10'b0100001001;
mem2[5230] = 10'b0100001010;
mem2[5231] = 10'b0100001010;
mem2[5232] = 10'b0100001010;
mem2[5233] = 10'b0100001010;
mem2[5234] = 10'b0100001010;
mem2[5235] = 10'b0100001010;
mem2[5236] = 10'b0100001010;
mem2[5237] = 10'b0100001010;
mem2[5238] = 10'b0100001010;
mem2[5239] = 10'b0100001010;
mem2[5240] = 10'b0100001010;
mem2[5241] = 10'b0100001011;
mem2[5242] = 10'b0100001011;
mem2[5243] = 10'b0100001011;
mem2[5244] = 10'b0100001011;
mem2[5245] = 10'b0100001011;
mem2[5246] = 10'b0100001011;
mem2[5247] = 10'b0100001011;
mem2[5248] = 10'b0100001011;
mem2[5249] = 10'b0100001011;
mem2[5250] = 10'b0100001011;
mem2[5251] = 10'b0100001100;
mem2[5252] = 10'b0100001100;
mem2[5253] = 10'b0100001100;
mem2[5254] = 10'b0100001100;
mem2[5255] = 10'b0100001100;
mem2[5256] = 10'b0100001100;
mem2[5257] = 10'b0100001100;
mem2[5258] = 10'b0100001100;
mem2[5259] = 10'b0100001100;
mem2[5260] = 10'b0100001100;
mem2[5261] = 10'b0100001100;
mem2[5262] = 10'b0100001101;
mem2[5263] = 10'b0100001101;
mem2[5264] = 10'b0100001101;
mem2[5265] = 10'b0100001101;
mem2[5266] = 10'b0100001101;
mem2[5267] = 10'b0100001101;
mem2[5268] = 10'b0100001101;
mem2[5269] = 10'b0100001101;
mem2[5270] = 10'b0100001101;
mem2[5271] = 10'b0100001101;
mem2[5272] = 10'b0100001101;
mem2[5273] = 10'b0100001110;
mem2[5274] = 10'b0100001110;
mem2[5275] = 10'b0100001110;
mem2[5276] = 10'b0100001110;
mem2[5277] = 10'b0100001110;
mem2[5278] = 10'b0100001110;
mem2[5279] = 10'b0100001110;
mem2[5280] = 10'b0100001110;
mem2[5281] = 10'b0100001110;
mem2[5282] = 10'b0100001110;
mem2[5283] = 10'b0100001110;
mem2[5284] = 10'b0100001111;
mem2[5285] = 10'b0100001111;
mem2[5286] = 10'b0100001111;
mem2[5287] = 10'b0100001111;
mem2[5288] = 10'b0100001111;
mem2[5289] = 10'b0100001111;
mem2[5290] = 10'b0100001111;
mem2[5291] = 10'b0100001111;
mem2[5292] = 10'b0100001111;
mem2[5293] = 10'b0100001111;
mem2[5294] = 10'b0100001111;
mem2[5295] = 10'b0100010000;
mem2[5296] = 10'b0100010000;
mem2[5297] = 10'b0100010000;
mem2[5298] = 10'b0100010000;
mem2[5299] = 10'b0100010000;
mem2[5300] = 10'b0100010000;
mem2[5301] = 10'b0100010000;
mem2[5302] = 10'b0100010000;
mem2[5303] = 10'b0100010000;
mem2[5304] = 10'b0100010000;
mem2[5305] = 10'b0100010000;
mem2[5306] = 10'b0100010001;
mem2[5307] = 10'b0100010001;
mem2[5308] = 10'b0100010001;
mem2[5309] = 10'b0100010001;
mem2[5310] = 10'b0100010001;
mem2[5311] = 10'b0100010001;
mem2[5312] = 10'b0100010001;
mem2[5313] = 10'b0100010001;
mem2[5314] = 10'b0100010001;
mem2[5315] = 10'b0100010001;
mem2[5316] = 10'b0100010010;
mem2[5317] = 10'b0100010010;
mem2[5318] = 10'b0100010010;
mem2[5319] = 10'b0100010010;
mem2[5320] = 10'b0100010010;
mem2[5321] = 10'b0100010010;
mem2[5322] = 10'b0100010010;
mem2[5323] = 10'b0100010010;
mem2[5324] = 10'b0100010010;
mem2[5325] = 10'b0100010010;
mem2[5326] = 10'b0100010010;
mem2[5327] = 10'b0100010011;
mem2[5328] = 10'b0100010011;
mem2[5329] = 10'b0100010011;
mem2[5330] = 10'b0100010011;
mem2[5331] = 10'b0100010011;
mem2[5332] = 10'b0100010011;
mem2[5333] = 10'b0100010011;
mem2[5334] = 10'b0100010011;
mem2[5335] = 10'b0100010011;
mem2[5336] = 10'b0100010011;
mem2[5337] = 10'b0100010011;
mem2[5338] = 10'b0100010100;
mem2[5339] = 10'b0100010100;
mem2[5340] = 10'b0100010100;
mem2[5341] = 10'b0100010100;
mem2[5342] = 10'b0100010100;
mem2[5343] = 10'b0100010100;
mem2[5344] = 10'b0100010100;
mem2[5345] = 10'b0100010100;
mem2[5346] = 10'b0100010100;
mem2[5347] = 10'b0100010100;
mem2[5348] = 10'b0100010100;
mem2[5349] = 10'b0100010101;
mem2[5350] = 10'b0100010101;
mem2[5351] = 10'b0100010101;
mem2[5352] = 10'b0100010101;
mem2[5353] = 10'b0100010101;
mem2[5354] = 10'b0100010101;
mem2[5355] = 10'b0100010101;
mem2[5356] = 10'b0100010101;
mem2[5357] = 10'b0100010101;
mem2[5358] = 10'b0100010101;
mem2[5359] = 10'b0100010110;
mem2[5360] = 10'b0100010110;
mem2[5361] = 10'b0100010110;
mem2[5362] = 10'b0100010110;
mem2[5363] = 10'b0100010110;
mem2[5364] = 10'b0100010110;
mem2[5365] = 10'b0100010110;
mem2[5366] = 10'b0100010110;
mem2[5367] = 10'b0100010110;
mem2[5368] = 10'b0100010110;
mem2[5369] = 10'b0100010110;
mem2[5370] = 10'b0100010111;
mem2[5371] = 10'b0100010111;
mem2[5372] = 10'b0100010111;
mem2[5373] = 10'b0100010111;
mem2[5374] = 10'b0100010111;
mem2[5375] = 10'b0100010111;
mem2[5376] = 10'b0100010111;
mem2[5377] = 10'b0100010111;
mem2[5378] = 10'b0100010111;
mem2[5379] = 10'b0100010111;
mem2[5380] = 10'b0100010111;
mem2[5381] = 10'b0100011000;
mem2[5382] = 10'b0100011000;
mem2[5383] = 10'b0100011000;
mem2[5384] = 10'b0100011000;
mem2[5385] = 10'b0100011000;
mem2[5386] = 10'b0100011000;
mem2[5387] = 10'b0100011000;
mem2[5388] = 10'b0100011000;
mem2[5389] = 10'b0100011000;
mem2[5390] = 10'b0100011000;
mem2[5391] = 10'b0100011000;
mem2[5392] = 10'b0100011001;
mem2[5393] = 10'b0100011001;
mem2[5394] = 10'b0100011001;
mem2[5395] = 10'b0100011001;
mem2[5396] = 10'b0100011001;
mem2[5397] = 10'b0100011001;
mem2[5398] = 10'b0100011001;
mem2[5399] = 10'b0100011001;
mem2[5400] = 10'b0100011001;
mem2[5401] = 10'b0100011001;
mem2[5402] = 10'b0100011010;
mem2[5403] = 10'b0100011010;
mem2[5404] = 10'b0100011010;
mem2[5405] = 10'b0100011010;
mem2[5406] = 10'b0100011010;
mem2[5407] = 10'b0100011010;
mem2[5408] = 10'b0100011010;
mem2[5409] = 10'b0100011010;
mem2[5410] = 10'b0100011010;
mem2[5411] = 10'b0100011010;
mem2[5412] = 10'b0100011010;
mem2[5413] = 10'b0100011011;
mem2[5414] = 10'b0100011011;
mem2[5415] = 10'b0100011011;
mem2[5416] = 10'b0100011011;
mem2[5417] = 10'b0100011011;
mem2[5418] = 10'b0100011011;
mem2[5419] = 10'b0100011011;
mem2[5420] = 10'b0100011011;
mem2[5421] = 10'b0100011011;
mem2[5422] = 10'b0100011011;
mem2[5423] = 10'b0100011011;
mem2[5424] = 10'b0100011100;
mem2[5425] = 10'b0100011100;
mem2[5426] = 10'b0100011100;
mem2[5427] = 10'b0100011100;
mem2[5428] = 10'b0100011100;
mem2[5429] = 10'b0100011100;
mem2[5430] = 10'b0100011100;
mem2[5431] = 10'b0100011100;
mem2[5432] = 10'b0100011100;
mem2[5433] = 10'b0100011100;
mem2[5434] = 10'b0100011101;
mem2[5435] = 10'b0100011101;
mem2[5436] = 10'b0100011101;
mem2[5437] = 10'b0100011101;
mem2[5438] = 10'b0100011101;
mem2[5439] = 10'b0100011101;
mem2[5440] = 10'b0100011101;
mem2[5441] = 10'b0100011101;
mem2[5442] = 10'b0100011101;
mem2[5443] = 10'b0100011101;
mem2[5444] = 10'b0100011101;
mem2[5445] = 10'b0100011110;
mem2[5446] = 10'b0100011110;
mem2[5447] = 10'b0100011110;
mem2[5448] = 10'b0100011110;
mem2[5449] = 10'b0100011110;
mem2[5450] = 10'b0100011110;
mem2[5451] = 10'b0100011110;
mem2[5452] = 10'b0100011110;
mem2[5453] = 10'b0100011110;
mem2[5454] = 10'b0100011110;
mem2[5455] = 10'b0100011110;
mem2[5456] = 10'b0100011111;
mem2[5457] = 10'b0100011111;
mem2[5458] = 10'b0100011111;
mem2[5459] = 10'b0100011111;
mem2[5460] = 10'b0100011111;
mem2[5461] = 10'b0100011111;
mem2[5462] = 10'b0100011111;
mem2[5463] = 10'b0100011111;
mem2[5464] = 10'b0100011111;
mem2[5465] = 10'b0100011111;
mem2[5466] = 10'b0100100000;
mem2[5467] = 10'b0100100000;
mem2[5468] = 10'b0100100000;
mem2[5469] = 10'b0100100000;
mem2[5470] = 10'b0100100000;
mem2[5471] = 10'b0100100000;
mem2[5472] = 10'b0100100000;
mem2[5473] = 10'b0100100000;
mem2[5474] = 10'b0100100000;
mem2[5475] = 10'b0100100000;
mem2[5476] = 10'b0100100000;
mem2[5477] = 10'b0100100001;
mem2[5478] = 10'b0100100001;
mem2[5479] = 10'b0100100001;
mem2[5480] = 10'b0100100001;
mem2[5481] = 10'b0100100001;
mem2[5482] = 10'b0100100001;
mem2[5483] = 10'b0100100001;
mem2[5484] = 10'b0100100001;
mem2[5485] = 10'b0100100001;
mem2[5486] = 10'b0100100001;
mem2[5487] = 10'b0100100010;
mem2[5488] = 10'b0100100010;
mem2[5489] = 10'b0100100010;
mem2[5490] = 10'b0100100010;
mem2[5491] = 10'b0100100010;
mem2[5492] = 10'b0100100010;
mem2[5493] = 10'b0100100010;
mem2[5494] = 10'b0100100010;
mem2[5495] = 10'b0100100010;
mem2[5496] = 10'b0100100010;
mem2[5497] = 10'b0100100010;
mem2[5498] = 10'b0100100011;
mem2[5499] = 10'b0100100011;
mem2[5500] = 10'b0100100011;
mem2[5501] = 10'b0100100011;
mem2[5502] = 10'b0100100011;
mem2[5503] = 10'b0100100011;
mem2[5504] = 10'b0100100011;
mem2[5505] = 10'b0100100011;
mem2[5506] = 10'b0100100011;
mem2[5507] = 10'b0100100011;
mem2[5508] = 10'b0100100011;
mem2[5509] = 10'b0100100100;
mem2[5510] = 10'b0100100100;
mem2[5511] = 10'b0100100100;
mem2[5512] = 10'b0100100100;
mem2[5513] = 10'b0100100100;
mem2[5514] = 10'b0100100100;
mem2[5515] = 10'b0100100100;
mem2[5516] = 10'b0100100100;
mem2[5517] = 10'b0100100100;
mem2[5518] = 10'b0100100100;
mem2[5519] = 10'b0100100101;
mem2[5520] = 10'b0100100101;
mem2[5521] = 10'b0100100101;
mem2[5522] = 10'b0100100101;
mem2[5523] = 10'b0100100101;
mem2[5524] = 10'b0100100101;
mem2[5525] = 10'b0100100101;
mem2[5526] = 10'b0100100101;
mem2[5527] = 10'b0100100101;
mem2[5528] = 10'b0100100101;
mem2[5529] = 10'b0100100101;
mem2[5530] = 10'b0100100110;
mem2[5531] = 10'b0100100110;
mem2[5532] = 10'b0100100110;
mem2[5533] = 10'b0100100110;
mem2[5534] = 10'b0100100110;
mem2[5535] = 10'b0100100110;
mem2[5536] = 10'b0100100110;
mem2[5537] = 10'b0100100110;
mem2[5538] = 10'b0100100110;
mem2[5539] = 10'b0100100110;
mem2[5540] = 10'b0100100111;
mem2[5541] = 10'b0100100111;
mem2[5542] = 10'b0100100111;
mem2[5543] = 10'b0100100111;
mem2[5544] = 10'b0100100111;
mem2[5545] = 10'b0100100111;
mem2[5546] = 10'b0100100111;
mem2[5547] = 10'b0100100111;
mem2[5548] = 10'b0100100111;
mem2[5549] = 10'b0100100111;
mem2[5550] = 10'b0100100111;
mem2[5551] = 10'b0100101000;
mem2[5552] = 10'b0100101000;
mem2[5553] = 10'b0100101000;
mem2[5554] = 10'b0100101000;
mem2[5555] = 10'b0100101000;
mem2[5556] = 10'b0100101000;
mem2[5557] = 10'b0100101000;
mem2[5558] = 10'b0100101000;
mem2[5559] = 10'b0100101000;
mem2[5560] = 10'b0100101000;
mem2[5561] = 10'b0100101001;
mem2[5562] = 10'b0100101001;
mem2[5563] = 10'b0100101001;
mem2[5564] = 10'b0100101001;
mem2[5565] = 10'b0100101001;
mem2[5566] = 10'b0100101001;
mem2[5567] = 10'b0100101001;
mem2[5568] = 10'b0100101001;
mem2[5569] = 10'b0100101001;
mem2[5570] = 10'b0100101001;
mem2[5571] = 10'b0100101001;
mem2[5572] = 10'b0100101010;
mem2[5573] = 10'b0100101010;
mem2[5574] = 10'b0100101010;
mem2[5575] = 10'b0100101010;
mem2[5576] = 10'b0100101010;
mem2[5577] = 10'b0100101010;
mem2[5578] = 10'b0100101010;
mem2[5579] = 10'b0100101010;
mem2[5580] = 10'b0100101010;
mem2[5581] = 10'b0100101010;
mem2[5582] = 10'b0100101011;
mem2[5583] = 10'b0100101011;
mem2[5584] = 10'b0100101011;
mem2[5585] = 10'b0100101011;
mem2[5586] = 10'b0100101011;
mem2[5587] = 10'b0100101011;
mem2[5588] = 10'b0100101011;
mem2[5589] = 10'b0100101011;
mem2[5590] = 10'b0100101011;
mem2[5591] = 10'b0100101011;
mem2[5592] = 10'b0100101011;
mem2[5593] = 10'b0100101100;
mem2[5594] = 10'b0100101100;
mem2[5595] = 10'b0100101100;
mem2[5596] = 10'b0100101100;
mem2[5597] = 10'b0100101100;
mem2[5598] = 10'b0100101100;
mem2[5599] = 10'b0100101100;
mem2[5600] = 10'b0100101100;
mem2[5601] = 10'b0100101100;
mem2[5602] = 10'b0100101100;
mem2[5603] = 10'b0100101101;
mem2[5604] = 10'b0100101101;
mem2[5605] = 10'b0100101101;
mem2[5606] = 10'b0100101101;
mem2[5607] = 10'b0100101101;
mem2[5608] = 10'b0100101101;
mem2[5609] = 10'b0100101101;
mem2[5610] = 10'b0100101101;
mem2[5611] = 10'b0100101101;
mem2[5612] = 10'b0100101101;
mem2[5613] = 10'b0100101101;
mem2[5614] = 10'b0100101110;
mem2[5615] = 10'b0100101110;
mem2[5616] = 10'b0100101110;
mem2[5617] = 10'b0100101110;
mem2[5618] = 10'b0100101110;
mem2[5619] = 10'b0100101110;
mem2[5620] = 10'b0100101110;
mem2[5621] = 10'b0100101110;
mem2[5622] = 10'b0100101110;
mem2[5623] = 10'b0100101110;
mem2[5624] = 10'b0100101111;
mem2[5625] = 10'b0100101111;
mem2[5626] = 10'b0100101111;
mem2[5627] = 10'b0100101111;
mem2[5628] = 10'b0100101111;
mem2[5629] = 10'b0100101111;
mem2[5630] = 10'b0100101111;
mem2[5631] = 10'b0100101111;
mem2[5632] = 10'b0100101111;
mem2[5633] = 10'b0100101111;
mem2[5634] = 10'b0100101111;
mem2[5635] = 10'b0100110000;
mem2[5636] = 10'b0100110000;
mem2[5637] = 10'b0100110000;
mem2[5638] = 10'b0100110000;
mem2[5639] = 10'b0100110000;
mem2[5640] = 10'b0100110000;
mem2[5641] = 10'b0100110000;
mem2[5642] = 10'b0100110000;
mem2[5643] = 10'b0100110000;
mem2[5644] = 10'b0100110000;
mem2[5645] = 10'b0100110001;
mem2[5646] = 10'b0100110001;
mem2[5647] = 10'b0100110001;
mem2[5648] = 10'b0100110001;
mem2[5649] = 10'b0100110001;
mem2[5650] = 10'b0100110001;
mem2[5651] = 10'b0100110001;
mem2[5652] = 10'b0100110001;
mem2[5653] = 10'b0100110001;
mem2[5654] = 10'b0100110001;
mem2[5655] = 10'b0100110001;
mem2[5656] = 10'b0100110010;
mem2[5657] = 10'b0100110010;
mem2[5658] = 10'b0100110010;
mem2[5659] = 10'b0100110010;
mem2[5660] = 10'b0100110010;
mem2[5661] = 10'b0100110010;
mem2[5662] = 10'b0100110010;
mem2[5663] = 10'b0100110010;
mem2[5664] = 10'b0100110010;
mem2[5665] = 10'b0100110010;
mem2[5666] = 10'b0100110011;
mem2[5667] = 10'b0100110011;
mem2[5668] = 10'b0100110011;
mem2[5669] = 10'b0100110011;
mem2[5670] = 10'b0100110011;
mem2[5671] = 10'b0100110011;
mem2[5672] = 10'b0100110011;
mem2[5673] = 10'b0100110011;
mem2[5674] = 10'b0100110011;
mem2[5675] = 10'b0100110011;
mem2[5676] = 10'b0100110100;
mem2[5677] = 10'b0100110100;
mem2[5678] = 10'b0100110100;
mem2[5679] = 10'b0100110100;
mem2[5680] = 10'b0100110100;
mem2[5681] = 10'b0100110100;
mem2[5682] = 10'b0100110100;
mem2[5683] = 10'b0100110100;
mem2[5684] = 10'b0100110100;
mem2[5685] = 10'b0100110100;
mem2[5686] = 10'b0100110100;
mem2[5687] = 10'b0100110101;
mem2[5688] = 10'b0100110101;
mem2[5689] = 10'b0100110101;
mem2[5690] = 10'b0100110101;
mem2[5691] = 10'b0100110101;
mem2[5692] = 10'b0100110101;
mem2[5693] = 10'b0100110101;
mem2[5694] = 10'b0100110101;
mem2[5695] = 10'b0100110101;
mem2[5696] = 10'b0100110101;
mem2[5697] = 10'b0100110110;
mem2[5698] = 10'b0100110110;
mem2[5699] = 10'b0100110110;
mem2[5700] = 10'b0100110110;
mem2[5701] = 10'b0100110110;
mem2[5702] = 10'b0100110110;
mem2[5703] = 10'b0100110110;
mem2[5704] = 10'b0100110110;
mem2[5705] = 10'b0100110110;
mem2[5706] = 10'b0100110110;
mem2[5707] = 10'b0100110110;
mem2[5708] = 10'b0100110111;
mem2[5709] = 10'b0100110111;
mem2[5710] = 10'b0100110111;
mem2[5711] = 10'b0100110111;
mem2[5712] = 10'b0100110111;
mem2[5713] = 10'b0100110111;
mem2[5714] = 10'b0100110111;
mem2[5715] = 10'b0100110111;
mem2[5716] = 10'b0100110111;
mem2[5717] = 10'b0100110111;
mem2[5718] = 10'b0100111000;
mem2[5719] = 10'b0100111000;
mem2[5720] = 10'b0100111000;
mem2[5721] = 10'b0100111000;
mem2[5722] = 10'b0100111000;
mem2[5723] = 10'b0100111000;
mem2[5724] = 10'b0100111000;
mem2[5725] = 10'b0100111000;
mem2[5726] = 10'b0100111000;
mem2[5727] = 10'b0100111000;
mem2[5728] = 10'b0100111001;
mem2[5729] = 10'b0100111001;
mem2[5730] = 10'b0100111001;
mem2[5731] = 10'b0100111001;
mem2[5732] = 10'b0100111001;
mem2[5733] = 10'b0100111001;
mem2[5734] = 10'b0100111001;
mem2[5735] = 10'b0100111001;
mem2[5736] = 10'b0100111001;
mem2[5737] = 10'b0100111001;
mem2[5738] = 10'b0100111001;
mem2[5739] = 10'b0100111010;
mem2[5740] = 10'b0100111010;
mem2[5741] = 10'b0100111010;
mem2[5742] = 10'b0100111010;
mem2[5743] = 10'b0100111010;
mem2[5744] = 10'b0100111010;
mem2[5745] = 10'b0100111010;
mem2[5746] = 10'b0100111010;
mem2[5747] = 10'b0100111010;
mem2[5748] = 10'b0100111010;
mem2[5749] = 10'b0100111011;
mem2[5750] = 10'b0100111011;
mem2[5751] = 10'b0100111011;
mem2[5752] = 10'b0100111011;
mem2[5753] = 10'b0100111011;
mem2[5754] = 10'b0100111011;
mem2[5755] = 10'b0100111011;
mem2[5756] = 10'b0100111011;
mem2[5757] = 10'b0100111011;
mem2[5758] = 10'b0100111011;
mem2[5759] = 10'b0100111100;
mem2[5760] = 10'b0100111100;
mem2[5761] = 10'b0100111100;
mem2[5762] = 10'b0100111100;
mem2[5763] = 10'b0100111100;
mem2[5764] = 10'b0100111100;
mem2[5765] = 10'b0100111100;
mem2[5766] = 10'b0100111100;
mem2[5767] = 10'b0100111100;
mem2[5768] = 10'b0100111100;
mem2[5769] = 10'b0100111100;
mem2[5770] = 10'b0100111101;
mem2[5771] = 10'b0100111101;
mem2[5772] = 10'b0100111101;
mem2[5773] = 10'b0100111101;
mem2[5774] = 10'b0100111101;
mem2[5775] = 10'b0100111101;
mem2[5776] = 10'b0100111101;
mem2[5777] = 10'b0100111101;
mem2[5778] = 10'b0100111101;
mem2[5779] = 10'b0100111101;
mem2[5780] = 10'b0100111110;
mem2[5781] = 10'b0100111110;
mem2[5782] = 10'b0100111110;
mem2[5783] = 10'b0100111110;
mem2[5784] = 10'b0100111110;
mem2[5785] = 10'b0100111110;
mem2[5786] = 10'b0100111110;
mem2[5787] = 10'b0100111110;
mem2[5788] = 10'b0100111110;
mem2[5789] = 10'b0100111110;
mem2[5790] = 10'b0100111111;
mem2[5791] = 10'b0100111111;
mem2[5792] = 10'b0100111111;
mem2[5793] = 10'b0100111111;
mem2[5794] = 10'b0100111111;
mem2[5795] = 10'b0100111111;
mem2[5796] = 10'b0100111111;
mem2[5797] = 10'b0100111111;
mem2[5798] = 10'b0100111111;
mem2[5799] = 10'b0100111111;
mem2[5800] = 10'b0100111111;
mem2[5801] = 10'b0101000000;
mem2[5802] = 10'b0101000000;
mem2[5803] = 10'b0101000000;
mem2[5804] = 10'b0101000000;
mem2[5805] = 10'b0101000000;
mem2[5806] = 10'b0101000000;
mem2[5807] = 10'b0101000000;
mem2[5808] = 10'b0101000000;
mem2[5809] = 10'b0101000000;
mem2[5810] = 10'b0101000000;
mem2[5811] = 10'b0101000001;
mem2[5812] = 10'b0101000001;
mem2[5813] = 10'b0101000001;
mem2[5814] = 10'b0101000001;
mem2[5815] = 10'b0101000001;
mem2[5816] = 10'b0101000001;
mem2[5817] = 10'b0101000001;
mem2[5818] = 10'b0101000001;
mem2[5819] = 10'b0101000001;
mem2[5820] = 10'b0101000001;
mem2[5821] = 10'b0101000010;
mem2[5822] = 10'b0101000010;
mem2[5823] = 10'b0101000010;
mem2[5824] = 10'b0101000010;
mem2[5825] = 10'b0101000010;
mem2[5826] = 10'b0101000010;
mem2[5827] = 10'b0101000010;
mem2[5828] = 10'b0101000010;
mem2[5829] = 10'b0101000010;
mem2[5830] = 10'b0101000010;
mem2[5831] = 10'b0101000010;
mem2[5832] = 10'b0101000011;
mem2[5833] = 10'b0101000011;
mem2[5834] = 10'b0101000011;
mem2[5835] = 10'b0101000011;
mem2[5836] = 10'b0101000011;
mem2[5837] = 10'b0101000011;
mem2[5838] = 10'b0101000011;
mem2[5839] = 10'b0101000011;
mem2[5840] = 10'b0101000011;
mem2[5841] = 10'b0101000011;
mem2[5842] = 10'b0101000100;
mem2[5843] = 10'b0101000100;
mem2[5844] = 10'b0101000100;
mem2[5845] = 10'b0101000100;
mem2[5846] = 10'b0101000100;
mem2[5847] = 10'b0101000100;
mem2[5848] = 10'b0101000100;
mem2[5849] = 10'b0101000100;
mem2[5850] = 10'b0101000100;
mem2[5851] = 10'b0101000100;
mem2[5852] = 10'b0101000101;
mem2[5853] = 10'b0101000101;
mem2[5854] = 10'b0101000101;
mem2[5855] = 10'b0101000101;
mem2[5856] = 10'b0101000101;
mem2[5857] = 10'b0101000101;
mem2[5858] = 10'b0101000101;
mem2[5859] = 10'b0101000101;
mem2[5860] = 10'b0101000101;
mem2[5861] = 10'b0101000101;
mem2[5862] = 10'b0101000110;
mem2[5863] = 10'b0101000110;
mem2[5864] = 10'b0101000110;
mem2[5865] = 10'b0101000110;
mem2[5866] = 10'b0101000110;
mem2[5867] = 10'b0101000110;
mem2[5868] = 10'b0101000110;
mem2[5869] = 10'b0101000110;
mem2[5870] = 10'b0101000110;
mem2[5871] = 10'b0101000110;
mem2[5872] = 10'b0101000110;
mem2[5873] = 10'b0101000111;
mem2[5874] = 10'b0101000111;
mem2[5875] = 10'b0101000111;
mem2[5876] = 10'b0101000111;
mem2[5877] = 10'b0101000111;
mem2[5878] = 10'b0101000111;
mem2[5879] = 10'b0101000111;
mem2[5880] = 10'b0101000111;
mem2[5881] = 10'b0101000111;
mem2[5882] = 10'b0101000111;
mem2[5883] = 10'b0101001000;
mem2[5884] = 10'b0101001000;
mem2[5885] = 10'b0101001000;
mem2[5886] = 10'b0101001000;
mem2[5887] = 10'b0101001000;
mem2[5888] = 10'b0101001000;
mem2[5889] = 10'b0101001000;
mem2[5890] = 10'b0101001000;
mem2[5891] = 10'b0101001000;
mem2[5892] = 10'b0101001000;
mem2[5893] = 10'b0101001001;
mem2[5894] = 10'b0101001001;
mem2[5895] = 10'b0101001001;
mem2[5896] = 10'b0101001001;
mem2[5897] = 10'b0101001001;
mem2[5898] = 10'b0101001001;
mem2[5899] = 10'b0101001001;
mem2[5900] = 10'b0101001001;
mem2[5901] = 10'b0101001001;
mem2[5902] = 10'b0101001001;
mem2[5903] = 10'b0101001010;
mem2[5904] = 10'b0101001010;
mem2[5905] = 10'b0101001010;
mem2[5906] = 10'b0101001010;
mem2[5907] = 10'b0101001010;
mem2[5908] = 10'b0101001010;
mem2[5909] = 10'b0101001010;
mem2[5910] = 10'b0101001010;
mem2[5911] = 10'b0101001010;
mem2[5912] = 10'b0101001010;
mem2[5913] = 10'b0101001011;
mem2[5914] = 10'b0101001011;
mem2[5915] = 10'b0101001011;
mem2[5916] = 10'b0101001011;
mem2[5917] = 10'b0101001011;
mem2[5918] = 10'b0101001011;
mem2[5919] = 10'b0101001011;
mem2[5920] = 10'b0101001011;
mem2[5921] = 10'b0101001011;
mem2[5922] = 10'b0101001011;
mem2[5923] = 10'b0101001011;
mem2[5924] = 10'b0101001100;
mem2[5925] = 10'b0101001100;
mem2[5926] = 10'b0101001100;
mem2[5927] = 10'b0101001100;
mem2[5928] = 10'b0101001100;
mem2[5929] = 10'b0101001100;
mem2[5930] = 10'b0101001100;
mem2[5931] = 10'b0101001100;
mem2[5932] = 10'b0101001100;
mem2[5933] = 10'b0101001100;
mem2[5934] = 10'b0101001101;
mem2[5935] = 10'b0101001101;
mem2[5936] = 10'b0101001101;
mem2[5937] = 10'b0101001101;
mem2[5938] = 10'b0101001101;
mem2[5939] = 10'b0101001101;
mem2[5940] = 10'b0101001101;
mem2[5941] = 10'b0101001101;
mem2[5942] = 10'b0101001101;
mem2[5943] = 10'b0101001101;
mem2[5944] = 10'b0101001110;
mem2[5945] = 10'b0101001110;
mem2[5946] = 10'b0101001110;
mem2[5947] = 10'b0101001110;
mem2[5948] = 10'b0101001110;
mem2[5949] = 10'b0101001110;
mem2[5950] = 10'b0101001110;
mem2[5951] = 10'b0101001110;
mem2[5952] = 10'b0101001110;
mem2[5953] = 10'b0101001110;
mem2[5954] = 10'b0101001111;
mem2[5955] = 10'b0101001111;
mem2[5956] = 10'b0101001111;
mem2[5957] = 10'b0101001111;
mem2[5958] = 10'b0101001111;
mem2[5959] = 10'b0101001111;
mem2[5960] = 10'b0101001111;
mem2[5961] = 10'b0101001111;
mem2[5962] = 10'b0101001111;
mem2[5963] = 10'b0101001111;
mem2[5964] = 10'b0101010000;
mem2[5965] = 10'b0101010000;
mem2[5966] = 10'b0101010000;
mem2[5967] = 10'b0101010000;
mem2[5968] = 10'b0101010000;
mem2[5969] = 10'b0101010000;
mem2[5970] = 10'b0101010000;
mem2[5971] = 10'b0101010000;
mem2[5972] = 10'b0101010000;
mem2[5973] = 10'b0101010000;
mem2[5974] = 10'b0101010000;
mem2[5975] = 10'b0101010001;
mem2[5976] = 10'b0101010001;
mem2[5977] = 10'b0101010001;
mem2[5978] = 10'b0101010001;
mem2[5979] = 10'b0101010001;
mem2[5980] = 10'b0101010001;
mem2[5981] = 10'b0101010001;
mem2[5982] = 10'b0101010001;
mem2[5983] = 10'b0101010001;
mem2[5984] = 10'b0101010001;
mem2[5985] = 10'b0101010010;
mem2[5986] = 10'b0101010010;
mem2[5987] = 10'b0101010010;
mem2[5988] = 10'b0101010010;
mem2[5989] = 10'b0101010010;
mem2[5990] = 10'b0101010010;
mem2[5991] = 10'b0101010010;
mem2[5992] = 10'b0101010010;
mem2[5993] = 10'b0101010010;
mem2[5994] = 10'b0101010010;
mem2[5995] = 10'b0101010011;
mem2[5996] = 10'b0101010011;
mem2[5997] = 10'b0101010011;
mem2[5998] = 10'b0101010011;
mem2[5999] = 10'b0101010011;
mem2[6000] = 10'b0101010011;
mem2[6001] = 10'b0101010011;
mem2[6002] = 10'b0101010011;
mem2[6003] = 10'b0101010011;
mem2[6004] = 10'b0101010011;
mem2[6005] = 10'b0101010100;
mem2[6006] = 10'b0101010100;
mem2[6007] = 10'b0101010100;
mem2[6008] = 10'b0101010100;
mem2[6009] = 10'b0101010100;
mem2[6010] = 10'b0101010100;
mem2[6011] = 10'b0101010100;
mem2[6012] = 10'b0101010100;
mem2[6013] = 10'b0101010100;
mem2[6014] = 10'b0101010100;
mem2[6015] = 10'b0101010101;
mem2[6016] = 10'b0101010101;
mem2[6017] = 10'b0101010101;
mem2[6018] = 10'b0101010101;
mem2[6019] = 10'b0101010101;
mem2[6020] = 10'b0101010101;
mem2[6021] = 10'b0101010101;
mem2[6022] = 10'b0101010101;
mem2[6023] = 10'b0101010101;
mem2[6024] = 10'b0101010101;
mem2[6025] = 10'b0101010110;
mem2[6026] = 10'b0101010110;
mem2[6027] = 10'b0101010110;
mem2[6028] = 10'b0101010110;
mem2[6029] = 10'b0101010110;
mem2[6030] = 10'b0101010110;
mem2[6031] = 10'b0101010110;
mem2[6032] = 10'b0101010110;
mem2[6033] = 10'b0101010110;
mem2[6034] = 10'b0101010110;
mem2[6035] = 10'b0101010111;
mem2[6036] = 10'b0101010111;
mem2[6037] = 10'b0101010111;
mem2[6038] = 10'b0101010111;
mem2[6039] = 10'b0101010111;
mem2[6040] = 10'b0101010111;
mem2[6041] = 10'b0101010111;
mem2[6042] = 10'b0101010111;
mem2[6043] = 10'b0101010111;
mem2[6044] = 10'b0101010111;
mem2[6045] = 10'b0101011000;
mem2[6046] = 10'b0101011000;
mem2[6047] = 10'b0101011000;
mem2[6048] = 10'b0101011000;
mem2[6049] = 10'b0101011000;
mem2[6050] = 10'b0101011000;
mem2[6051] = 10'b0101011000;
mem2[6052] = 10'b0101011000;
mem2[6053] = 10'b0101011000;
mem2[6054] = 10'b0101011000;
mem2[6055] = 10'b0101011000;
mem2[6056] = 10'b0101011001;
mem2[6057] = 10'b0101011001;
mem2[6058] = 10'b0101011001;
mem2[6059] = 10'b0101011001;
mem2[6060] = 10'b0101011001;
mem2[6061] = 10'b0101011001;
mem2[6062] = 10'b0101011001;
mem2[6063] = 10'b0101011001;
mem2[6064] = 10'b0101011001;
mem2[6065] = 10'b0101011001;
mem2[6066] = 10'b0101011010;
mem2[6067] = 10'b0101011010;
mem2[6068] = 10'b0101011010;
mem2[6069] = 10'b0101011010;
mem2[6070] = 10'b0101011010;
mem2[6071] = 10'b0101011010;
mem2[6072] = 10'b0101011010;
mem2[6073] = 10'b0101011010;
mem2[6074] = 10'b0101011010;
mem2[6075] = 10'b0101011010;
mem2[6076] = 10'b0101011011;
mem2[6077] = 10'b0101011011;
mem2[6078] = 10'b0101011011;
mem2[6079] = 10'b0101011011;
mem2[6080] = 10'b0101011011;
mem2[6081] = 10'b0101011011;
mem2[6082] = 10'b0101011011;
mem2[6083] = 10'b0101011011;
mem2[6084] = 10'b0101011011;
mem2[6085] = 10'b0101011011;
mem2[6086] = 10'b0101011100;
mem2[6087] = 10'b0101011100;
mem2[6088] = 10'b0101011100;
mem2[6089] = 10'b0101011100;
mem2[6090] = 10'b0101011100;
mem2[6091] = 10'b0101011100;
mem2[6092] = 10'b0101011100;
mem2[6093] = 10'b0101011100;
mem2[6094] = 10'b0101011100;
mem2[6095] = 10'b0101011100;
mem2[6096] = 10'b0101011101;
mem2[6097] = 10'b0101011101;
mem2[6098] = 10'b0101011101;
mem2[6099] = 10'b0101011101;
mem2[6100] = 10'b0101011101;
mem2[6101] = 10'b0101011101;
mem2[6102] = 10'b0101011101;
mem2[6103] = 10'b0101011101;
mem2[6104] = 10'b0101011101;
mem2[6105] = 10'b0101011101;
mem2[6106] = 10'b0101011110;
mem2[6107] = 10'b0101011110;
mem2[6108] = 10'b0101011110;
mem2[6109] = 10'b0101011110;
mem2[6110] = 10'b0101011110;
mem2[6111] = 10'b0101011110;
mem2[6112] = 10'b0101011110;
mem2[6113] = 10'b0101011110;
mem2[6114] = 10'b0101011110;
mem2[6115] = 10'b0101011110;
mem2[6116] = 10'b0101011111;
mem2[6117] = 10'b0101011111;
mem2[6118] = 10'b0101011111;
mem2[6119] = 10'b0101011111;
mem2[6120] = 10'b0101011111;
mem2[6121] = 10'b0101011111;
mem2[6122] = 10'b0101011111;
mem2[6123] = 10'b0101011111;
mem2[6124] = 10'b0101011111;
mem2[6125] = 10'b0101011111;
mem2[6126] = 10'b0101100000;
mem2[6127] = 10'b0101100000;
mem2[6128] = 10'b0101100000;
mem2[6129] = 10'b0101100000;
mem2[6130] = 10'b0101100000;
mem2[6131] = 10'b0101100000;
mem2[6132] = 10'b0101100000;
mem2[6133] = 10'b0101100000;
mem2[6134] = 10'b0101100000;
mem2[6135] = 10'b0101100000;
mem2[6136] = 10'b0101100001;
mem2[6137] = 10'b0101100001;
mem2[6138] = 10'b0101100001;
mem2[6139] = 10'b0101100001;
mem2[6140] = 10'b0101100001;
mem2[6141] = 10'b0101100001;
mem2[6142] = 10'b0101100001;
mem2[6143] = 10'b0101100001;
mem2[6144] = 10'b0101100001;
mem2[6145] = 10'b0101100001;
mem2[6146] = 10'b0101100010;
mem2[6147] = 10'b0101100010;
mem2[6148] = 10'b0101100010;
mem2[6149] = 10'b0101100010;
mem2[6150] = 10'b0101100010;
mem2[6151] = 10'b0101100010;
mem2[6152] = 10'b0101100010;
mem2[6153] = 10'b0101100010;
mem2[6154] = 10'b0101100010;
mem2[6155] = 10'b0101100010;
mem2[6156] = 10'b0101100011;
mem2[6157] = 10'b0101100011;
mem2[6158] = 10'b0101100011;
mem2[6159] = 10'b0101100011;
mem2[6160] = 10'b0101100011;
mem2[6161] = 10'b0101100011;
mem2[6162] = 10'b0101100011;
mem2[6163] = 10'b0101100011;
mem2[6164] = 10'b0101100011;
mem2[6165] = 10'b0101100011;
mem2[6166] = 10'b0101100100;
mem2[6167] = 10'b0101100100;
mem2[6168] = 10'b0101100100;
mem2[6169] = 10'b0101100100;
mem2[6170] = 10'b0101100100;
mem2[6171] = 10'b0101100100;
mem2[6172] = 10'b0101100100;
mem2[6173] = 10'b0101100100;
mem2[6174] = 10'b0101100100;
mem2[6175] = 10'b0101100100;
mem2[6176] = 10'b0101100101;
mem2[6177] = 10'b0101100101;
mem2[6178] = 10'b0101100101;
mem2[6179] = 10'b0101100101;
mem2[6180] = 10'b0101100101;
mem2[6181] = 10'b0101100101;
mem2[6182] = 10'b0101100101;
mem2[6183] = 10'b0101100101;
mem2[6184] = 10'b0101100101;
mem2[6185] = 10'b0101100101;
mem2[6186] = 10'b0101100110;
mem2[6187] = 10'b0101100110;
mem2[6188] = 10'b0101100110;
mem2[6189] = 10'b0101100110;
mem2[6190] = 10'b0101100110;
mem2[6191] = 10'b0101100110;
mem2[6192] = 10'b0101100110;
mem2[6193] = 10'b0101100110;
mem2[6194] = 10'b0101100110;
mem2[6195] = 10'b0101100110;
mem2[6196] = 10'b0101100111;
mem2[6197] = 10'b0101100111;
mem2[6198] = 10'b0101100111;
mem2[6199] = 10'b0101100111;
mem2[6200] = 10'b0101100111;
mem2[6201] = 10'b0101100111;
mem2[6202] = 10'b0101100111;
mem2[6203] = 10'b0101100111;
mem2[6204] = 10'b0101100111;
mem2[6205] = 10'b0101100111;
mem2[6206] = 10'b0101101000;
mem2[6207] = 10'b0101101000;
mem2[6208] = 10'b0101101000;
mem2[6209] = 10'b0101101000;
mem2[6210] = 10'b0101101000;
mem2[6211] = 10'b0101101000;
mem2[6212] = 10'b0101101000;
mem2[6213] = 10'b0101101000;
mem2[6214] = 10'b0101101000;
mem2[6215] = 10'b0101101000;
mem2[6216] = 10'b0101101001;
mem2[6217] = 10'b0101101001;
mem2[6218] = 10'b0101101001;
mem2[6219] = 10'b0101101001;
mem2[6220] = 10'b0101101001;
mem2[6221] = 10'b0101101001;
mem2[6222] = 10'b0101101001;
mem2[6223] = 10'b0101101001;
mem2[6224] = 10'b0101101001;
mem2[6225] = 10'b0101101001;
mem2[6226] = 10'b0101101010;
mem2[6227] = 10'b0101101010;
mem2[6228] = 10'b0101101010;
mem2[6229] = 10'b0101101010;
mem2[6230] = 10'b0101101010;
mem2[6231] = 10'b0101101010;
mem2[6232] = 10'b0101101010;
mem2[6233] = 10'b0101101010;
mem2[6234] = 10'b0101101010;
mem2[6235] = 10'b0101101010;
mem2[6236] = 10'b0101101011;
mem2[6237] = 10'b0101101011;
mem2[6238] = 10'b0101101011;
mem2[6239] = 10'b0101101011;
mem2[6240] = 10'b0101101011;
mem2[6241] = 10'b0101101011;
mem2[6242] = 10'b0101101011;
mem2[6243] = 10'b0101101011;
mem2[6244] = 10'b0101101011;
mem2[6245] = 10'b0101101011;
mem2[6246] = 10'b0101101100;
mem2[6247] = 10'b0101101100;
mem2[6248] = 10'b0101101100;
mem2[6249] = 10'b0101101100;
mem2[6250] = 10'b0101101100;
mem2[6251] = 10'b0101101100;
mem2[6252] = 10'b0101101100;
mem2[6253] = 10'b0101101100;
mem2[6254] = 10'b0101101100;
mem2[6255] = 10'b0101101100;
mem2[6256] = 10'b0101101101;
mem2[6257] = 10'b0101101101;
mem2[6258] = 10'b0101101101;
mem2[6259] = 10'b0101101101;
mem2[6260] = 10'b0101101101;
mem2[6261] = 10'b0101101101;
mem2[6262] = 10'b0101101101;
mem2[6263] = 10'b0101101101;
mem2[6264] = 10'b0101101101;
mem2[6265] = 10'b0101101101;
mem2[6266] = 10'b0101101110;
mem2[6267] = 10'b0101101110;
mem2[6268] = 10'b0101101110;
mem2[6269] = 10'b0101101110;
mem2[6270] = 10'b0101101110;
mem2[6271] = 10'b0101101110;
mem2[6272] = 10'b0101101110;
mem2[6273] = 10'b0101101110;
mem2[6274] = 10'b0101101110;
mem2[6275] = 10'b0101101110;
mem2[6276] = 10'b0101101111;
mem2[6277] = 10'b0101101111;
mem2[6278] = 10'b0101101111;
mem2[6279] = 10'b0101101111;
mem2[6280] = 10'b0101101111;
mem2[6281] = 10'b0101101111;
mem2[6282] = 10'b0101101111;
mem2[6283] = 10'b0101101111;
mem2[6284] = 10'b0101101111;
mem2[6285] = 10'b0101101111;
mem2[6286] = 10'b0101110000;
mem2[6287] = 10'b0101110000;
mem2[6288] = 10'b0101110000;
mem2[6289] = 10'b0101110000;
mem2[6290] = 10'b0101110000;
mem2[6291] = 10'b0101110000;
mem2[6292] = 10'b0101110000;
mem2[6293] = 10'b0101110000;
mem2[6294] = 10'b0101110000;
mem2[6295] = 10'b0101110000;
mem2[6296] = 10'b0101110001;
mem2[6297] = 10'b0101110001;
mem2[6298] = 10'b0101110001;
mem2[6299] = 10'b0101110001;
mem2[6300] = 10'b0101110001;
mem2[6301] = 10'b0101110001;
mem2[6302] = 10'b0101110001;
mem2[6303] = 10'b0101110001;
mem2[6304] = 10'b0101110001;
mem2[6305] = 10'b0101110001;
mem2[6306] = 10'b0101110010;
mem2[6307] = 10'b0101110010;
mem2[6308] = 10'b0101110010;
mem2[6309] = 10'b0101110010;
mem2[6310] = 10'b0101110010;
mem2[6311] = 10'b0101110010;
mem2[6312] = 10'b0101110010;
mem2[6313] = 10'b0101110010;
mem2[6314] = 10'b0101110010;
mem2[6315] = 10'b0101110010;
mem2[6316] = 10'b0101110011;
mem2[6317] = 10'b0101110011;
mem2[6318] = 10'b0101110011;
mem2[6319] = 10'b0101110011;
mem2[6320] = 10'b0101110011;
mem2[6321] = 10'b0101110011;
mem2[6322] = 10'b0101110011;
mem2[6323] = 10'b0101110011;
mem2[6324] = 10'b0101110011;
mem2[6325] = 10'b0101110011;
mem2[6326] = 10'b0101110100;
mem2[6327] = 10'b0101110100;
mem2[6328] = 10'b0101110100;
mem2[6329] = 10'b0101110100;
mem2[6330] = 10'b0101110100;
mem2[6331] = 10'b0101110100;
mem2[6332] = 10'b0101110100;
mem2[6333] = 10'b0101110100;
mem2[6334] = 10'b0101110100;
mem2[6335] = 10'b0101110100;
mem2[6336] = 10'b0101110101;
mem2[6337] = 10'b0101110101;
mem2[6338] = 10'b0101110101;
mem2[6339] = 10'b0101110101;
mem2[6340] = 10'b0101110101;
mem2[6341] = 10'b0101110101;
mem2[6342] = 10'b0101110101;
mem2[6343] = 10'b0101110101;
mem2[6344] = 10'b0101110101;
mem2[6345] = 10'b0101110101;
mem2[6346] = 10'b0101110110;
mem2[6347] = 10'b0101110110;
mem2[6348] = 10'b0101110110;
mem2[6349] = 10'b0101110110;
mem2[6350] = 10'b0101110110;
mem2[6351] = 10'b0101110110;
mem2[6352] = 10'b0101110110;
mem2[6353] = 10'b0101110110;
mem2[6354] = 10'b0101110110;
mem2[6355] = 10'b0101110110;
mem2[6356] = 10'b0101110111;
mem2[6357] = 10'b0101110111;
mem2[6358] = 10'b0101110111;
mem2[6359] = 10'b0101110111;
mem2[6360] = 10'b0101110111;
mem2[6361] = 10'b0101110111;
mem2[6362] = 10'b0101110111;
mem2[6363] = 10'b0101110111;
mem2[6364] = 10'b0101110111;
mem2[6365] = 10'b0101110111;
mem2[6366] = 10'b0101111000;
mem2[6367] = 10'b0101111000;
mem2[6368] = 10'b0101111000;
mem2[6369] = 10'b0101111000;
mem2[6370] = 10'b0101111000;
mem2[6371] = 10'b0101111000;
mem2[6372] = 10'b0101111000;
mem2[6373] = 10'b0101111000;
mem2[6374] = 10'b0101111000;
mem2[6375] = 10'b0101111001;
mem2[6376] = 10'b0101111001;
mem2[6377] = 10'b0101111001;
mem2[6378] = 10'b0101111001;
mem2[6379] = 10'b0101111001;
mem2[6380] = 10'b0101111001;
mem2[6381] = 10'b0101111001;
mem2[6382] = 10'b0101111001;
mem2[6383] = 10'b0101111001;
mem2[6384] = 10'b0101111001;
mem2[6385] = 10'b0101111010;
mem2[6386] = 10'b0101111010;
mem2[6387] = 10'b0101111010;
mem2[6388] = 10'b0101111010;
mem2[6389] = 10'b0101111010;
mem2[6390] = 10'b0101111010;
mem2[6391] = 10'b0101111010;
mem2[6392] = 10'b0101111010;
mem2[6393] = 10'b0101111010;
mem2[6394] = 10'b0101111010;
mem2[6395] = 10'b0101111011;
mem2[6396] = 10'b0101111011;
mem2[6397] = 10'b0101111011;
mem2[6398] = 10'b0101111011;
mem2[6399] = 10'b0101111011;
mem2[6400] = 10'b0101111011;
mem2[6401] = 10'b0101111011;
mem2[6402] = 10'b0101111011;
mem2[6403] = 10'b0101111011;
mem2[6404] = 10'b0101111011;
mem2[6405] = 10'b0101111100;
mem2[6406] = 10'b0101111100;
mem2[6407] = 10'b0101111100;
mem2[6408] = 10'b0101111100;
mem2[6409] = 10'b0101111100;
mem2[6410] = 10'b0101111100;
mem2[6411] = 10'b0101111100;
mem2[6412] = 10'b0101111100;
mem2[6413] = 10'b0101111100;
mem2[6414] = 10'b0101111100;
mem2[6415] = 10'b0101111101;
mem2[6416] = 10'b0101111101;
mem2[6417] = 10'b0101111101;
mem2[6418] = 10'b0101111101;
mem2[6419] = 10'b0101111101;
mem2[6420] = 10'b0101111101;
mem2[6421] = 10'b0101111101;
mem2[6422] = 10'b0101111101;
mem2[6423] = 10'b0101111101;
mem2[6424] = 10'b0101111101;
mem2[6425] = 10'b0101111110;
mem2[6426] = 10'b0101111110;
mem2[6427] = 10'b0101111110;
mem2[6428] = 10'b0101111110;
mem2[6429] = 10'b0101111110;
mem2[6430] = 10'b0101111110;
mem2[6431] = 10'b0101111110;
mem2[6432] = 10'b0101111110;
mem2[6433] = 10'b0101111110;
mem2[6434] = 10'b0101111110;
mem2[6435] = 10'b0101111111;
mem2[6436] = 10'b0101111111;
mem2[6437] = 10'b0101111111;
mem2[6438] = 10'b0101111111;
mem2[6439] = 10'b0101111111;
mem2[6440] = 10'b0101111111;
mem2[6441] = 10'b0101111111;
mem2[6442] = 10'b0101111111;
mem2[6443] = 10'b0101111111;
mem2[6444] = 10'b0101111111;
mem2[6445] = 10'b0110000000;
mem2[6446] = 10'b0110000000;
mem2[6447] = 10'b0110000000;
mem2[6448] = 10'b0110000000;
mem2[6449] = 10'b0110000000;
mem2[6450] = 10'b0110000000;
mem2[6451] = 10'b0110000000;
mem2[6452] = 10'b0110000000;
mem2[6453] = 10'b0110000000;
mem2[6454] = 10'b0110000001;
mem2[6455] = 10'b0110000001;
mem2[6456] = 10'b0110000001;
mem2[6457] = 10'b0110000001;
mem2[6458] = 10'b0110000001;
mem2[6459] = 10'b0110000001;
mem2[6460] = 10'b0110000001;
mem2[6461] = 10'b0110000001;
mem2[6462] = 10'b0110000001;
mem2[6463] = 10'b0110000001;
mem2[6464] = 10'b0110000010;
mem2[6465] = 10'b0110000010;
mem2[6466] = 10'b0110000010;
mem2[6467] = 10'b0110000010;
mem2[6468] = 10'b0110000010;
mem2[6469] = 10'b0110000010;
mem2[6470] = 10'b0110000010;
mem2[6471] = 10'b0110000010;
mem2[6472] = 10'b0110000010;
mem2[6473] = 10'b0110000010;
mem2[6474] = 10'b0110000011;
mem2[6475] = 10'b0110000011;
mem2[6476] = 10'b0110000011;
mem2[6477] = 10'b0110000011;
mem2[6478] = 10'b0110000011;
mem2[6479] = 10'b0110000011;
mem2[6480] = 10'b0110000011;
mem2[6481] = 10'b0110000011;
mem2[6482] = 10'b0110000011;
mem2[6483] = 10'b0110000011;
mem2[6484] = 10'b0110000100;
mem2[6485] = 10'b0110000100;
mem2[6486] = 10'b0110000100;
mem2[6487] = 10'b0110000100;
mem2[6488] = 10'b0110000100;
mem2[6489] = 10'b0110000100;
mem2[6490] = 10'b0110000100;
mem2[6491] = 10'b0110000100;
mem2[6492] = 10'b0110000100;
mem2[6493] = 10'b0110000100;
mem2[6494] = 10'b0110000101;
mem2[6495] = 10'b0110000101;
mem2[6496] = 10'b0110000101;
mem2[6497] = 10'b0110000101;
mem2[6498] = 10'b0110000101;
mem2[6499] = 10'b0110000101;
mem2[6500] = 10'b0110000101;
mem2[6501] = 10'b0110000101;
mem2[6502] = 10'b0110000101;
mem2[6503] = 10'b0110000101;
mem2[6504] = 10'b0110000110;
mem2[6505] = 10'b0110000110;
mem2[6506] = 10'b0110000110;
mem2[6507] = 10'b0110000110;
mem2[6508] = 10'b0110000110;
mem2[6509] = 10'b0110000110;
mem2[6510] = 10'b0110000110;
mem2[6511] = 10'b0110000110;
mem2[6512] = 10'b0110000110;
mem2[6513] = 10'b0110000110;
mem2[6514] = 10'b0110000111;
mem2[6515] = 10'b0110000111;
mem2[6516] = 10'b0110000111;
mem2[6517] = 10'b0110000111;
mem2[6518] = 10'b0110000111;
mem2[6519] = 10'b0110000111;
mem2[6520] = 10'b0110000111;
mem2[6521] = 10'b0110000111;
mem2[6522] = 10'b0110000111;
mem2[6523] = 10'b0110001000;
mem2[6524] = 10'b0110001000;
mem2[6525] = 10'b0110001000;
mem2[6526] = 10'b0110001000;
mem2[6527] = 10'b0110001000;
mem2[6528] = 10'b0110001000;
mem2[6529] = 10'b0110001000;
mem2[6530] = 10'b0110001000;
mem2[6531] = 10'b0110001000;
mem2[6532] = 10'b0110001000;
mem2[6533] = 10'b0110001001;
mem2[6534] = 10'b0110001001;
mem2[6535] = 10'b0110001001;
mem2[6536] = 10'b0110001001;
mem2[6537] = 10'b0110001001;
mem2[6538] = 10'b0110001001;
mem2[6539] = 10'b0110001001;
mem2[6540] = 10'b0110001001;
mem2[6541] = 10'b0110001001;
mem2[6542] = 10'b0110001001;
mem2[6543] = 10'b0110001010;
mem2[6544] = 10'b0110001010;
mem2[6545] = 10'b0110001010;
mem2[6546] = 10'b0110001010;
mem2[6547] = 10'b0110001010;
mem2[6548] = 10'b0110001010;
mem2[6549] = 10'b0110001010;
mem2[6550] = 10'b0110001010;
mem2[6551] = 10'b0110001010;
mem2[6552] = 10'b0110001010;
mem2[6553] = 10'b0110001011;
mem2[6554] = 10'b0110001011;
mem2[6555] = 10'b0110001011;
mem2[6556] = 10'b0110001011;
mem2[6557] = 10'b0110001011;
mem2[6558] = 10'b0110001011;
mem2[6559] = 10'b0110001011;
mem2[6560] = 10'b0110001011;
mem2[6561] = 10'b0110001011;
mem2[6562] = 10'b0110001011;
mem2[6563] = 10'b0110001100;
mem2[6564] = 10'b0110001100;
mem2[6565] = 10'b0110001100;
mem2[6566] = 10'b0110001100;
mem2[6567] = 10'b0110001100;
mem2[6568] = 10'b0110001100;
mem2[6569] = 10'b0110001100;
mem2[6570] = 10'b0110001100;
mem2[6571] = 10'b0110001100;
mem2[6572] = 10'b0110001101;
mem2[6573] = 10'b0110001101;
mem2[6574] = 10'b0110001101;
mem2[6575] = 10'b0110001101;
mem2[6576] = 10'b0110001101;
mem2[6577] = 10'b0110001101;
mem2[6578] = 10'b0110001101;
mem2[6579] = 10'b0110001101;
mem2[6580] = 10'b0110001101;
mem2[6581] = 10'b0110001101;
mem2[6582] = 10'b0110001110;
mem2[6583] = 10'b0110001110;
mem2[6584] = 10'b0110001110;
mem2[6585] = 10'b0110001110;
mem2[6586] = 10'b0110001110;
mem2[6587] = 10'b0110001110;
mem2[6588] = 10'b0110001110;
mem2[6589] = 10'b0110001110;
mem2[6590] = 10'b0110001110;
mem2[6591] = 10'b0110001110;
mem2[6592] = 10'b0110001111;
mem2[6593] = 10'b0110001111;
mem2[6594] = 10'b0110001111;
mem2[6595] = 10'b0110001111;
mem2[6596] = 10'b0110001111;
mem2[6597] = 10'b0110001111;
mem2[6598] = 10'b0110001111;
mem2[6599] = 10'b0110001111;
mem2[6600] = 10'b0110001111;
mem2[6601] = 10'b0110001111;
mem2[6602] = 10'b0110010000;
mem2[6603] = 10'b0110010000;
mem2[6604] = 10'b0110010000;
mem2[6605] = 10'b0110010000;
mem2[6606] = 10'b0110010000;
mem2[6607] = 10'b0110010000;
mem2[6608] = 10'b0110010000;
mem2[6609] = 10'b0110010000;
mem2[6610] = 10'b0110010000;
mem2[6611] = 10'b0110010000;
mem2[6612] = 10'b0110010001;
mem2[6613] = 10'b0110010001;
mem2[6614] = 10'b0110010001;
mem2[6615] = 10'b0110010001;
mem2[6616] = 10'b0110010001;
mem2[6617] = 10'b0110010001;
mem2[6618] = 10'b0110010001;
mem2[6619] = 10'b0110010001;
mem2[6620] = 10'b0110010001;
mem2[6621] = 10'b0110010010;
mem2[6622] = 10'b0110010010;
mem2[6623] = 10'b0110010010;
mem2[6624] = 10'b0110010010;
mem2[6625] = 10'b0110010010;
mem2[6626] = 10'b0110010010;
mem2[6627] = 10'b0110010010;
mem2[6628] = 10'b0110010010;
mem2[6629] = 10'b0110010010;
mem2[6630] = 10'b0110010010;
mem2[6631] = 10'b0110010011;
mem2[6632] = 10'b0110010011;
mem2[6633] = 10'b0110010011;
mem2[6634] = 10'b0110010011;
mem2[6635] = 10'b0110010011;
mem2[6636] = 10'b0110010011;
mem2[6637] = 10'b0110010011;
mem2[6638] = 10'b0110010011;
mem2[6639] = 10'b0110010011;
mem2[6640] = 10'b0110010011;
mem2[6641] = 10'b0110010100;
mem2[6642] = 10'b0110010100;
mem2[6643] = 10'b0110010100;
mem2[6644] = 10'b0110010100;
mem2[6645] = 10'b0110010100;
mem2[6646] = 10'b0110010100;
mem2[6647] = 10'b0110010100;
mem2[6648] = 10'b0110010100;
mem2[6649] = 10'b0110010100;
mem2[6650] = 10'b0110010100;
mem2[6651] = 10'b0110010101;
mem2[6652] = 10'b0110010101;
mem2[6653] = 10'b0110010101;
mem2[6654] = 10'b0110010101;
mem2[6655] = 10'b0110010101;
mem2[6656] = 10'b0110010101;
mem2[6657] = 10'b0110010101;
mem2[6658] = 10'b0110010101;
mem2[6659] = 10'b0110010101;
mem2[6660] = 10'b0110010110;
mem2[6661] = 10'b0110010110;
mem2[6662] = 10'b0110010110;
mem2[6663] = 10'b0110010110;
mem2[6664] = 10'b0110010110;
mem2[6665] = 10'b0110010110;
mem2[6666] = 10'b0110010110;
mem2[6667] = 10'b0110010110;
mem2[6668] = 10'b0110010110;
mem2[6669] = 10'b0110010110;
mem2[6670] = 10'b0110010111;
mem2[6671] = 10'b0110010111;
mem2[6672] = 10'b0110010111;
mem2[6673] = 10'b0110010111;
mem2[6674] = 10'b0110010111;
mem2[6675] = 10'b0110010111;
mem2[6676] = 10'b0110010111;
mem2[6677] = 10'b0110010111;
mem2[6678] = 10'b0110010111;
mem2[6679] = 10'b0110010111;
mem2[6680] = 10'b0110011000;
mem2[6681] = 10'b0110011000;
mem2[6682] = 10'b0110011000;
mem2[6683] = 10'b0110011000;
mem2[6684] = 10'b0110011000;
mem2[6685] = 10'b0110011000;
mem2[6686] = 10'b0110011000;
mem2[6687] = 10'b0110011000;
mem2[6688] = 10'b0110011000;
mem2[6689] = 10'b0110011000;
mem2[6690] = 10'b0110011001;
mem2[6691] = 10'b0110011001;
mem2[6692] = 10'b0110011001;
mem2[6693] = 10'b0110011001;
mem2[6694] = 10'b0110011001;
mem2[6695] = 10'b0110011001;
mem2[6696] = 10'b0110011001;
mem2[6697] = 10'b0110011001;
mem2[6698] = 10'b0110011001;
mem2[6699] = 10'b0110011010;
mem2[6700] = 10'b0110011010;
mem2[6701] = 10'b0110011010;
mem2[6702] = 10'b0110011010;
mem2[6703] = 10'b0110011010;
mem2[6704] = 10'b0110011010;
mem2[6705] = 10'b0110011010;
mem2[6706] = 10'b0110011010;
mem2[6707] = 10'b0110011010;
mem2[6708] = 10'b0110011010;
mem2[6709] = 10'b0110011011;
mem2[6710] = 10'b0110011011;
mem2[6711] = 10'b0110011011;
mem2[6712] = 10'b0110011011;
mem2[6713] = 10'b0110011011;
mem2[6714] = 10'b0110011011;
mem2[6715] = 10'b0110011011;
mem2[6716] = 10'b0110011011;
mem2[6717] = 10'b0110011011;
mem2[6718] = 10'b0110011011;
mem2[6719] = 10'b0110011100;
mem2[6720] = 10'b0110011100;
mem2[6721] = 10'b0110011100;
mem2[6722] = 10'b0110011100;
mem2[6723] = 10'b0110011100;
mem2[6724] = 10'b0110011100;
mem2[6725] = 10'b0110011100;
mem2[6726] = 10'b0110011100;
mem2[6727] = 10'b0110011100;
mem2[6728] = 10'b0110011100;
mem2[6729] = 10'b0110011101;
mem2[6730] = 10'b0110011101;
mem2[6731] = 10'b0110011101;
mem2[6732] = 10'b0110011101;
mem2[6733] = 10'b0110011101;
mem2[6734] = 10'b0110011101;
mem2[6735] = 10'b0110011101;
mem2[6736] = 10'b0110011101;
mem2[6737] = 10'b0110011101;
mem2[6738] = 10'b0110011110;
mem2[6739] = 10'b0110011110;
mem2[6740] = 10'b0110011110;
mem2[6741] = 10'b0110011110;
mem2[6742] = 10'b0110011110;
mem2[6743] = 10'b0110011110;
mem2[6744] = 10'b0110011110;
mem2[6745] = 10'b0110011110;
mem2[6746] = 10'b0110011110;
mem2[6747] = 10'b0110011110;
mem2[6748] = 10'b0110011111;
mem2[6749] = 10'b0110011111;
mem2[6750] = 10'b0110011111;
mem2[6751] = 10'b0110011111;
mem2[6752] = 10'b0110011111;
mem2[6753] = 10'b0110011111;
mem2[6754] = 10'b0110011111;
mem2[6755] = 10'b0110011111;
mem2[6756] = 10'b0110011111;
mem2[6757] = 10'b0110011111;
mem2[6758] = 10'b0110100000;
mem2[6759] = 10'b0110100000;
mem2[6760] = 10'b0110100000;
mem2[6761] = 10'b0110100000;
mem2[6762] = 10'b0110100000;
mem2[6763] = 10'b0110100000;
mem2[6764] = 10'b0110100000;
mem2[6765] = 10'b0110100000;
mem2[6766] = 10'b0110100000;
mem2[6767] = 10'b0110100000;
mem2[6768] = 10'b0110100001;
mem2[6769] = 10'b0110100001;
mem2[6770] = 10'b0110100001;
mem2[6771] = 10'b0110100001;
mem2[6772] = 10'b0110100001;
mem2[6773] = 10'b0110100001;
mem2[6774] = 10'b0110100001;
mem2[6775] = 10'b0110100001;
mem2[6776] = 10'b0110100001;
mem2[6777] = 10'b0110100010;
mem2[6778] = 10'b0110100010;
mem2[6779] = 10'b0110100010;
mem2[6780] = 10'b0110100010;
mem2[6781] = 10'b0110100010;
mem2[6782] = 10'b0110100010;
mem2[6783] = 10'b0110100010;
mem2[6784] = 10'b0110100010;
mem2[6785] = 10'b0110100010;
mem2[6786] = 10'b0110100010;
mem2[6787] = 10'b0110100011;
mem2[6788] = 10'b0110100011;
mem2[6789] = 10'b0110100011;
mem2[6790] = 10'b0110100011;
mem2[6791] = 10'b0110100011;
mem2[6792] = 10'b0110100011;
mem2[6793] = 10'b0110100011;
mem2[6794] = 10'b0110100011;
mem2[6795] = 10'b0110100011;
mem2[6796] = 10'b0110100011;
mem2[6797] = 10'b0110100100;
mem2[6798] = 10'b0110100100;
mem2[6799] = 10'b0110100100;
mem2[6800] = 10'b0110100100;
mem2[6801] = 10'b0110100100;
mem2[6802] = 10'b0110100100;
mem2[6803] = 10'b0110100100;
mem2[6804] = 10'b0110100100;
mem2[6805] = 10'b0110100100;
mem2[6806] = 10'b0110100101;
mem2[6807] = 10'b0110100101;
mem2[6808] = 10'b0110100101;
mem2[6809] = 10'b0110100101;
mem2[6810] = 10'b0110100101;
mem2[6811] = 10'b0110100101;
mem2[6812] = 10'b0110100101;
mem2[6813] = 10'b0110100101;
mem2[6814] = 10'b0110100101;
mem2[6815] = 10'b0110100101;
mem2[6816] = 10'b0110100110;
mem2[6817] = 10'b0110100110;
mem2[6818] = 10'b0110100110;
mem2[6819] = 10'b0110100110;
mem2[6820] = 10'b0110100110;
mem2[6821] = 10'b0110100110;
mem2[6822] = 10'b0110100110;
mem2[6823] = 10'b0110100110;
mem2[6824] = 10'b0110100110;
mem2[6825] = 10'b0110100110;
mem2[6826] = 10'b0110100111;
mem2[6827] = 10'b0110100111;
mem2[6828] = 10'b0110100111;
mem2[6829] = 10'b0110100111;
mem2[6830] = 10'b0110100111;
mem2[6831] = 10'b0110100111;
mem2[6832] = 10'b0110100111;
mem2[6833] = 10'b0110100111;
mem2[6834] = 10'b0110100111;
mem2[6835] = 10'b0110101000;
mem2[6836] = 10'b0110101000;
mem2[6837] = 10'b0110101000;
mem2[6838] = 10'b0110101000;
mem2[6839] = 10'b0110101000;
mem2[6840] = 10'b0110101000;
mem2[6841] = 10'b0110101000;
mem2[6842] = 10'b0110101000;
mem2[6843] = 10'b0110101000;
mem2[6844] = 10'b0110101000;
mem2[6845] = 10'b0110101001;
mem2[6846] = 10'b0110101001;
mem2[6847] = 10'b0110101001;
mem2[6848] = 10'b0110101001;
mem2[6849] = 10'b0110101001;
mem2[6850] = 10'b0110101001;
mem2[6851] = 10'b0110101001;
mem2[6852] = 10'b0110101001;
mem2[6853] = 10'b0110101001;
mem2[6854] = 10'b0110101001;
mem2[6855] = 10'b0110101010;
mem2[6856] = 10'b0110101010;
mem2[6857] = 10'b0110101010;
mem2[6858] = 10'b0110101010;
mem2[6859] = 10'b0110101010;
mem2[6860] = 10'b0110101010;
mem2[6861] = 10'b0110101010;
mem2[6862] = 10'b0110101010;
mem2[6863] = 10'b0110101010;
mem2[6864] = 10'b0110101010;
mem2[6865] = 10'b0110101011;
mem2[6866] = 10'b0110101011;
mem2[6867] = 10'b0110101011;
mem2[6868] = 10'b0110101011;
mem2[6869] = 10'b0110101011;
mem2[6870] = 10'b0110101011;
mem2[6871] = 10'b0110101011;
mem2[6872] = 10'b0110101011;
mem2[6873] = 10'b0110101011;
mem2[6874] = 10'b0110101100;
mem2[6875] = 10'b0110101100;
mem2[6876] = 10'b0110101100;
mem2[6877] = 10'b0110101100;
mem2[6878] = 10'b0110101100;
mem2[6879] = 10'b0110101100;
mem2[6880] = 10'b0110101100;
mem2[6881] = 10'b0110101100;
mem2[6882] = 10'b0110101100;
mem2[6883] = 10'b0110101100;
mem2[6884] = 10'b0110101101;
mem2[6885] = 10'b0110101101;
mem2[6886] = 10'b0110101101;
mem2[6887] = 10'b0110101101;
mem2[6888] = 10'b0110101101;
mem2[6889] = 10'b0110101101;
mem2[6890] = 10'b0110101101;
mem2[6891] = 10'b0110101101;
mem2[6892] = 10'b0110101101;
mem2[6893] = 10'b0110101101;
mem2[6894] = 10'b0110101110;
mem2[6895] = 10'b0110101110;
mem2[6896] = 10'b0110101110;
mem2[6897] = 10'b0110101110;
mem2[6898] = 10'b0110101110;
mem2[6899] = 10'b0110101110;
mem2[6900] = 10'b0110101110;
mem2[6901] = 10'b0110101110;
mem2[6902] = 10'b0110101110;
mem2[6903] = 10'b0110101111;
mem2[6904] = 10'b0110101111;
mem2[6905] = 10'b0110101111;
mem2[6906] = 10'b0110101111;
mem2[6907] = 10'b0110101111;
mem2[6908] = 10'b0110101111;
mem2[6909] = 10'b0110101111;
mem2[6910] = 10'b0110101111;
mem2[6911] = 10'b0110101111;
mem2[6912] = 10'b0110101111;
mem2[6913] = 10'b0110110000;
mem2[6914] = 10'b0110110000;
mem2[6915] = 10'b0110110000;
mem2[6916] = 10'b0110110000;
mem2[6917] = 10'b0110110000;
mem2[6918] = 10'b0110110000;
mem2[6919] = 10'b0110110000;
mem2[6920] = 10'b0110110000;
mem2[6921] = 10'b0110110000;
mem2[6922] = 10'b0110110000;
mem2[6923] = 10'b0110110001;
mem2[6924] = 10'b0110110001;
mem2[6925] = 10'b0110110001;
mem2[6926] = 10'b0110110001;
mem2[6927] = 10'b0110110001;
mem2[6928] = 10'b0110110001;
mem2[6929] = 10'b0110110001;
mem2[6930] = 10'b0110110001;
mem2[6931] = 10'b0110110001;
mem2[6932] = 10'b0110110010;
mem2[6933] = 10'b0110110010;
mem2[6934] = 10'b0110110010;
mem2[6935] = 10'b0110110010;
mem2[6936] = 10'b0110110010;
mem2[6937] = 10'b0110110010;
mem2[6938] = 10'b0110110010;
mem2[6939] = 10'b0110110010;
mem2[6940] = 10'b0110110010;
mem2[6941] = 10'b0110110010;
mem2[6942] = 10'b0110110011;
mem2[6943] = 10'b0110110011;
mem2[6944] = 10'b0110110011;
mem2[6945] = 10'b0110110011;
mem2[6946] = 10'b0110110011;
mem2[6947] = 10'b0110110011;
mem2[6948] = 10'b0110110011;
mem2[6949] = 10'b0110110011;
mem2[6950] = 10'b0110110011;
mem2[6951] = 10'b0110110011;
mem2[6952] = 10'b0110110100;
mem2[6953] = 10'b0110110100;
mem2[6954] = 10'b0110110100;
mem2[6955] = 10'b0110110100;
mem2[6956] = 10'b0110110100;
mem2[6957] = 10'b0110110100;
mem2[6958] = 10'b0110110100;
mem2[6959] = 10'b0110110100;
mem2[6960] = 10'b0110110100;
mem2[6961] = 10'b0110110101;
mem2[6962] = 10'b0110110101;
mem2[6963] = 10'b0110110101;
mem2[6964] = 10'b0110110101;
mem2[6965] = 10'b0110110101;
mem2[6966] = 10'b0110110101;
mem2[6967] = 10'b0110110101;
mem2[6968] = 10'b0110110101;
mem2[6969] = 10'b0110110101;
mem2[6970] = 10'b0110110101;
mem2[6971] = 10'b0110110110;
mem2[6972] = 10'b0110110110;
mem2[6973] = 10'b0110110110;
mem2[6974] = 10'b0110110110;
mem2[6975] = 10'b0110110110;
mem2[6976] = 10'b0110110110;
mem2[6977] = 10'b0110110110;
mem2[6978] = 10'b0110110110;
mem2[6979] = 10'b0110110110;
mem2[6980] = 10'b0110110110;
mem2[6981] = 10'b0110110111;
mem2[6982] = 10'b0110110111;
mem2[6983] = 10'b0110110111;
mem2[6984] = 10'b0110110111;
mem2[6985] = 10'b0110110111;
mem2[6986] = 10'b0110110111;
mem2[6987] = 10'b0110110111;
mem2[6988] = 10'b0110110111;
mem2[6989] = 10'b0110110111;
mem2[6990] = 10'b0110111000;
mem2[6991] = 10'b0110111000;
mem2[6992] = 10'b0110111000;
mem2[6993] = 10'b0110111000;
mem2[6994] = 10'b0110111000;
mem2[6995] = 10'b0110111000;
mem2[6996] = 10'b0110111000;
mem2[6997] = 10'b0110111000;
mem2[6998] = 10'b0110111000;
mem2[6999] = 10'b0110111000;
mem2[7000] = 10'b0110111001;
mem2[7001] = 10'b0110111001;
mem2[7002] = 10'b0110111001;
mem2[7003] = 10'b0110111001;
mem2[7004] = 10'b0110111001;
mem2[7005] = 10'b0110111001;
mem2[7006] = 10'b0110111001;
mem2[7007] = 10'b0110111001;
mem2[7008] = 10'b0110111001;
mem2[7009] = 10'b0110111010;
mem2[7010] = 10'b0110111010;
mem2[7011] = 10'b0110111010;
mem2[7012] = 10'b0110111010;
mem2[7013] = 10'b0110111010;
mem2[7014] = 10'b0110111010;
mem2[7015] = 10'b0110111010;
mem2[7016] = 10'b0110111010;
mem2[7017] = 10'b0110111010;
mem2[7018] = 10'b0110111010;
mem2[7019] = 10'b0110111011;
mem2[7020] = 10'b0110111011;
mem2[7021] = 10'b0110111011;
mem2[7022] = 10'b0110111011;
mem2[7023] = 10'b0110111011;
mem2[7024] = 10'b0110111011;
mem2[7025] = 10'b0110111011;
mem2[7026] = 10'b0110111011;
mem2[7027] = 10'b0110111011;
mem2[7028] = 10'b0110111011;
mem2[7029] = 10'b0110111100;
mem2[7030] = 10'b0110111100;
mem2[7031] = 10'b0110111100;
mem2[7032] = 10'b0110111100;
mem2[7033] = 10'b0110111100;
mem2[7034] = 10'b0110111100;
mem2[7035] = 10'b0110111100;
mem2[7036] = 10'b0110111100;
mem2[7037] = 10'b0110111100;
mem2[7038] = 10'b0110111101;
mem2[7039] = 10'b0110111101;
mem2[7040] = 10'b0110111101;
mem2[7041] = 10'b0110111101;
mem2[7042] = 10'b0110111101;
mem2[7043] = 10'b0110111101;
mem2[7044] = 10'b0110111101;
mem2[7045] = 10'b0110111101;
mem2[7046] = 10'b0110111101;
mem2[7047] = 10'b0110111101;
mem2[7048] = 10'b0110111110;
mem2[7049] = 10'b0110111110;
mem2[7050] = 10'b0110111110;
mem2[7051] = 10'b0110111110;
mem2[7052] = 10'b0110111110;
mem2[7053] = 10'b0110111110;
mem2[7054] = 10'b0110111110;
mem2[7055] = 10'b0110111110;
mem2[7056] = 10'b0110111110;
mem2[7057] = 10'b0110111110;
mem2[7058] = 10'b0110111111;
mem2[7059] = 10'b0110111111;
mem2[7060] = 10'b0110111111;
mem2[7061] = 10'b0110111111;
mem2[7062] = 10'b0110111111;
mem2[7063] = 10'b0110111111;
mem2[7064] = 10'b0110111111;
mem2[7065] = 10'b0110111111;
mem2[7066] = 10'b0110111111;
mem2[7067] = 10'b0111000000;
mem2[7068] = 10'b0111000000;
mem2[7069] = 10'b0111000000;
mem2[7070] = 10'b0111000000;
mem2[7071] = 10'b0111000000;
mem2[7072] = 10'b0111000000;
mem2[7073] = 10'b0111000000;
mem2[7074] = 10'b0111000000;
mem2[7075] = 10'b0111000000;
mem2[7076] = 10'b0111000000;
mem2[7077] = 10'b0111000001;
mem2[7078] = 10'b0111000001;
mem2[7079] = 10'b0111000001;
mem2[7080] = 10'b0111000001;
mem2[7081] = 10'b0111000001;
mem2[7082] = 10'b0111000001;
mem2[7083] = 10'b0111000001;
mem2[7084] = 10'b0111000001;
mem2[7085] = 10'b0111000001;
mem2[7086] = 10'b0111000001;
mem2[7087] = 10'b0111000010;
mem2[7088] = 10'b0111000010;
mem2[7089] = 10'b0111000010;
mem2[7090] = 10'b0111000010;
mem2[7091] = 10'b0111000010;
mem2[7092] = 10'b0111000010;
mem2[7093] = 10'b0111000010;
mem2[7094] = 10'b0111000010;
mem2[7095] = 10'b0111000010;
mem2[7096] = 10'b0111000011;
mem2[7097] = 10'b0111000011;
mem2[7098] = 10'b0111000011;
mem2[7099] = 10'b0111000011;
mem2[7100] = 10'b0111000011;
mem2[7101] = 10'b0111000011;
mem2[7102] = 10'b0111000011;
mem2[7103] = 10'b0111000011;
mem2[7104] = 10'b0111000011;
mem2[7105] = 10'b0111000011;
mem2[7106] = 10'b0111000100;
mem2[7107] = 10'b0111000100;
mem2[7108] = 10'b0111000100;
mem2[7109] = 10'b0111000100;
mem2[7110] = 10'b0111000100;
mem2[7111] = 10'b0111000100;
mem2[7112] = 10'b0111000100;
mem2[7113] = 10'b0111000100;
mem2[7114] = 10'b0111000100;
mem2[7115] = 10'b0111000101;
mem2[7116] = 10'b0111000101;
mem2[7117] = 10'b0111000101;
mem2[7118] = 10'b0111000101;
mem2[7119] = 10'b0111000101;
mem2[7120] = 10'b0111000101;
mem2[7121] = 10'b0111000101;
mem2[7122] = 10'b0111000101;
mem2[7123] = 10'b0111000101;
mem2[7124] = 10'b0111000101;
mem2[7125] = 10'b0111000110;
mem2[7126] = 10'b0111000110;
mem2[7127] = 10'b0111000110;
mem2[7128] = 10'b0111000110;
mem2[7129] = 10'b0111000110;
mem2[7130] = 10'b0111000110;
mem2[7131] = 10'b0111000110;
mem2[7132] = 10'b0111000110;
mem2[7133] = 10'b0111000110;
mem2[7134] = 10'b0111000110;
mem2[7135] = 10'b0111000111;
mem2[7136] = 10'b0111000111;
mem2[7137] = 10'b0111000111;
mem2[7138] = 10'b0111000111;
mem2[7139] = 10'b0111000111;
mem2[7140] = 10'b0111000111;
mem2[7141] = 10'b0111000111;
mem2[7142] = 10'b0111000111;
mem2[7143] = 10'b0111000111;
mem2[7144] = 10'b0111001000;
mem2[7145] = 10'b0111001000;
mem2[7146] = 10'b0111001000;
mem2[7147] = 10'b0111001000;
mem2[7148] = 10'b0111001000;
mem2[7149] = 10'b0111001000;
mem2[7150] = 10'b0111001000;
mem2[7151] = 10'b0111001000;
mem2[7152] = 10'b0111001000;
mem2[7153] = 10'b0111001000;
mem2[7154] = 10'b0111001001;
mem2[7155] = 10'b0111001001;
mem2[7156] = 10'b0111001001;
mem2[7157] = 10'b0111001001;
mem2[7158] = 10'b0111001001;
mem2[7159] = 10'b0111001001;
mem2[7160] = 10'b0111001001;
mem2[7161] = 10'b0111001001;
mem2[7162] = 10'b0111001001;
mem2[7163] = 10'b0111001010;
mem2[7164] = 10'b0111001010;
mem2[7165] = 10'b0111001010;
mem2[7166] = 10'b0111001010;
mem2[7167] = 10'b0111001010;
mem2[7168] = 10'b0111001010;
mem2[7169] = 10'b0111001010;
mem2[7170] = 10'b0111001010;
mem2[7171] = 10'b0111001010;
mem2[7172] = 10'b0111001010;
mem2[7173] = 10'b0111001011;
mem2[7174] = 10'b0111001011;
mem2[7175] = 10'b0111001011;
mem2[7176] = 10'b0111001011;
mem2[7177] = 10'b0111001011;
mem2[7178] = 10'b0111001011;
mem2[7179] = 10'b0111001011;
mem2[7180] = 10'b0111001011;
mem2[7181] = 10'b0111001011;
mem2[7182] = 10'b0111001011;
mem2[7183] = 10'b0111001100;
mem2[7184] = 10'b0111001100;
mem2[7185] = 10'b0111001100;
mem2[7186] = 10'b0111001100;
mem2[7187] = 10'b0111001100;
mem2[7188] = 10'b0111001100;
mem2[7189] = 10'b0111001100;
mem2[7190] = 10'b0111001100;
mem2[7191] = 10'b0111001100;
mem2[7192] = 10'b0111001101;
mem2[7193] = 10'b0111001101;
mem2[7194] = 10'b0111001101;
mem2[7195] = 10'b0111001101;
mem2[7196] = 10'b0111001101;
mem2[7197] = 10'b0111001101;
mem2[7198] = 10'b0111001101;
mem2[7199] = 10'b0111001101;
mem2[7200] = 10'b0111001101;
mem2[7201] = 10'b0111001101;
mem2[7202] = 10'b0111001110;
mem2[7203] = 10'b0111001110;
mem2[7204] = 10'b0111001110;
mem2[7205] = 10'b0111001110;
mem2[7206] = 10'b0111001110;
mem2[7207] = 10'b0111001110;
mem2[7208] = 10'b0111001110;
mem2[7209] = 10'b0111001110;
mem2[7210] = 10'b0111001110;
mem2[7211] = 10'b0111001111;
mem2[7212] = 10'b0111001111;
mem2[7213] = 10'b0111001111;
mem2[7214] = 10'b0111001111;
mem2[7215] = 10'b0111001111;
mem2[7216] = 10'b0111001111;
mem2[7217] = 10'b0111001111;
mem2[7218] = 10'b0111001111;
mem2[7219] = 10'b0111001111;
mem2[7220] = 10'b0111001111;
mem2[7221] = 10'b0111010000;
mem2[7222] = 10'b0111010000;
mem2[7223] = 10'b0111010000;
mem2[7224] = 10'b0111010000;
mem2[7225] = 10'b0111010000;
mem2[7226] = 10'b0111010000;
mem2[7227] = 10'b0111010000;
mem2[7228] = 10'b0111010000;
mem2[7229] = 10'b0111010000;
mem2[7230] = 10'b0111010000;
mem2[7231] = 10'b0111010001;
mem2[7232] = 10'b0111010001;
mem2[7233] = 10'b0111010001;
mem2[7234] = 10'b0111010001;
mem2[7235] = 10'b0111010001;
mem2[7236] = 10'b0111010001;
mem2[7237] = 10'b0111010001;
mem2[7238] = 10'b0111010001;
mem2[7239] = 10'b0111010001;
mem2[7240] = 10'b0111010010;
mem2[7241] = 10'b0111010010;
mem2[7242] = 10'b0111010010;
mem2[7243] = 10'b0111010010;
mem2[7244] = 10'b0111010010;
mem2[7245] = 10'b0111010010;
mem2[7246] = 10'b0111010010;
mem2[7247] = 10'b0111010010;
mem2[7248] = 10'b0111010010;
mem2[7249] = 10'b0111010010;
mem2[7250] = 10'b0111010011;
mem2[7251] = 10'b0111010011;
mem2[7252] = 10'b0111010011;
mem2[7253] = 10'b0111010011;
mem2[7254] = 10'b0111010011;
mem2[7255] = 10'b0111010011;
mem2[7256] = 10'b0111010011;
mem2[7257] = 10'b0111010011;
mem2[7258] = 10'b0111010011;
mem2[7259] = 10'b0111010100;
mem2[7260] = 10'b0111010100;
mem2[7261] = 10'b0111010100;
mem2[7262] = 10'b0111010100;
mem2[7263] = 10'b0111010100;
mem2[7264] = 10'b0111010100;
mem2[7265] = 10'b0111010100;
mem2[7266] = 10'b0111010100;
mem2[7267] = 10'b0111010100;
mem2[7268] = 10'b0111010100;
mem2[7269] = 10'b0111010101;
mem2[7270] = 10'b0111010101;
mem2[7271] = 10'b0111010101;
mem2[7272] = 10'b0111010101;
mem2[7273] = 10'b0111010101;
mem2[7274] = 10'b0111010101;
mem2[7275] = 10'b0111010101;
mem2[7276] = 10'b0111010101;
mem2[7277] = 10'b0111010101;
mem2[7278] = 10'b0111010110;
mem2[7279] = 10'b0111010110;
mem2[7280] = 10'b0111010110;
mem2[7281] = 10'b0111010110;
mem2[7282] = 10'b0111010110;
mem2[7283] = 10'b0111010110;
mem2[7284] = 10'b0111010110;
mem2[7285] = 10'b0111010110;
mem2[7286] = 10'b0111010110;
mem2[7287] = 10'b0111010110;
mem2[7288] = 10'b0111010111;
mem2[7289] = 10'b0111010111;
mem2[7290] = 10'b0111010111;
mem2[7291] = 10'b0111010111;
mem2[7292] = 10'b0111010111;
mem2[7293] = 10'b0111010111;
mem2[7294] = 10'b0111010111;
mem2[7295] = 10'b0111010111;
mem2[7296] = 10'b0111010111;
mem2[7297] = 10'b0111010111;
mem2[7298] = 10'b0111011000;
mem2[7299] = 10'b0111011000;
mem2[7300] = 10'b0111011000;
mem2[7301] = 10'b0111011000;
mem2[7302] = 10'b0111011000;
mem2[7303] = 10'b0111011000;
mem2[7304] = 10'b0111011000;
mem2[7305] = 10'b0111011000;
mem2[7306] = 10'b0111011000;
mem2[7307] = 10'b0111011001;
mem2[7308] = 10'b0111011001;
mem2[7309] = 10'b0111011001;
mem2[7310] = 10'b0111011001;
mem2[7311] = 10'b0111011001;
mem2[7312] = 10'b0111011001;
mem2[7313] = 10'b0111011001;
mem2[7314] = 10'b0111011001;
mem2[7315] = 10'b0111011001;
mem2[7316] = 10'b0111011001;
mem2[7317] = 10'b0111011010;
mem2[7318] = 10'b0111011010;
mem2[7319] = 10'b0111011010;
mem2[7320] = 10'b0111011010;
mem2[7321] = 10'b0111011010;
mem2[7322] = 10'b0111011010;
mem2[7323] = 10'b0111011010;
mem2[7324] = 10'b0111011010;
mem2[7325] = 10'b0111011010;
mem2[7326] = 10'b0111011011;
mem2[7327] = 10'b0111011011;
mem2[7328] = 10'b0111011011;
mem2[7329] = 10'b0111011011;
mem2[7330] = 10'b0111011011;
mem2[7331] = 10'b0111011011;
mem2[7332] = 10'b0111011011;
mem2[7333] = 10'b0111011011;
mem2[7334] = 10'b0111011011;
mem2[7335] = 10'b0111011011;
mem2[7336] = 10'b0111011100;
mem2[7337] = 10'b0111011100;
mem2[7338] = 10'b0111011100;
mem2[7339] = 10'b0111011100;
mem2[7340] = 10'b0111011100;
mem2[7341] = 10'b0111011100;
mem2[7342] = 10'b0111011100;
mem2[7343] = 10'b0111011100;
mem2[7344] = 10'b0111011100;
mem2[7345] = 10'b0111011100;
mem2[7346] = 10'b0111011101;
mem2[7347] = 10'b0111011101;
mem2[7348] = 10'b0111011101;
mem2[7349] = 10'b0111011101;
mem2[7350] = 10'b0111011101;
mem2[7351] = 10'b0111011101;
mem2[7352] = 10'b0111011101;
mem2[7353] = 10'b0111011101;
mem2[7354] = 10'b0111011101;
mem2[7355] = 10'b0111011110;
mem2[7356] = 10'b0111011110;
mem2[7357] = 10'b0111011110;
mem2[7358] = 10'b0111011110;
mem2[7359] = 10'b0111011110;
mem2[7360] = 10'b0111011110;
mem2[7361] = 10'b0111011110;
mem2[7362] = 10'b0111011110;
mem2[7363] = 10'b0111011110;
mem2[7364] = 10'b0111011110;
mem2[7365] = 10'b0111011111;
mem2[7366] = 10'b0111011111;
mem2[7367] = 10'b0111011111;
mem2[7368] = 10'b0111011111;
mem2[7369] = 10'b0111011111;
mem2[7370] = 10'b0111011111;
mem2[7371] = 10'b0111011111;
mem2[7372] = 10'b0111011111;
mem2[7373] = 10'b0111011111;
mem2[7374] = 10'b0111100000;
mem2[7375] = 10'b0111100000;
mem2[7376] = 10'b0111100000;
mem2[7377] = 10'b0111100000;
mem2[7378] = 10'b0111100000;
mem2[7379] = 10'b0111100000;
mem2[7380] = 10'b0111100000;
mem2[7381] = 10'b0111100000;
mem2[7382] = 10'b0111100000;
mem2[7383] = 10'b0111100000;
mem2[7384] = 10'b0111100001;
mem2[7385] = 10'b0111100001;
mem2[7386] = 10'b0111100001;
mem2[7387] = 10'b0111100001;
mem2[7388] = 10'b0111100001;
mem2[7389] = 10'b0111100001;
mem2[7390] = 10'b0111100001;
mem2[7391] = 10'b0111100001;
mem2[7392] = 10'b0111100001;
mem2[7393] = 10'b0111100010;
mem2[7394] = 10'b0111100010;
mem2[7395] = 10'b0111100010;
mem2[7396] = 10'b0111100010;
mem2[7397] = 10'b0111100010;
mem2[7398] = 10'b0111100010;
mem2[7399] = 10'b0111100010;
mem2[7400] = 10'b0111100010;
mem2[7401] = 10'b0111100010;
mem2[7402] = 10'b0111100010;
mem2[7403] = 10'b0111100011;
mem2[7404] = 10'b0111100011;
mem2[7405] = 10'b0111100011;
mem2[7406] = 10'b0111100011;
mem2[7407] = 10'b0111100011;
mem2[7408] = 10'b0111100011;
mem2[7409] = 10'b0111100011;
mem2[7410] = 10'b0111100011;
mem2[7411] = 10'b0111100011;
mem2[7412] = 10'b0111100100;
mem2[7413] = 10'b0111100100;
mem2[7414] = 10'b0111100100;
mem2[7415] = 10'b0111100100;
mem2[7416] = 10'b0111100100;
mem2[7417] = 10'b0111100100;
mem2[7418] = 10'b0111100100;
mem2[7419] = 10'b0111100100;
mem2[7420] = 10'b0111100100;
mem2[7421] = 10'b0111100100;
mem2[7422] = 10'b0111100101;
mem2[7423] = 10'b0111100101;
mem2[7424] = 10'b0111100101;
mem2[7425] = 10'b0111100101;
mem2[7426] = 10'b0111100101;
mem2[7427] = 10'b0111100101;
mem2[7428] = 10'b0111100101;
mem2[7429] = 10'b0111100101;
mem2[7430] = 10'b0111100101;
mem2[7431] = 10'b0111100101;
mem2[7432] = 10'b0111100110;
mem2[7433] = 10'b0111100110;
mem2[7434] = 10'b0111100110;
mem2[7435] = 10'b0111100110;
mem2[7436] = 10'b0111100110;
mem2[7437] = 10'b0111100110;
mem2[7438] = 10'b0111100110;
mem2[7439] = 10'b0111100110;
mem2[7440] = 10'b0111100110;
mem2[7441] = 10'b0111100111;
mem2[7442] = 10'b0111100111;
mem2[7443] = 10'b0111100111;
mem2[7444] = 10'b0111100111;
mem2[7445] = 10'b0111100111;
mem2[7446] = 10'b0111100111;
mem2[7447] = 10'b0111100111;
mem2[7448] = 10'b0111100111;
mem2[7449] = 10'b0111100111;
mem2[7450] = 10'b0111100111;
mem2[7451] = 10'b0111101000;
mem2[7452] = 10'b0111101000;
mem2[7453] = 10'b0111101000;
mem2[7454] = 10'b0111101000;
mem2[7455] = 10'b0111101000;
mem2[7456] = 10'b0111101000;
mem2[7457] = 10'b0111101000;
mem2[7458] = 10'b0111101000;
mem2[7459] = 10'b0111101000;
mem2[7460] = 10'b0111101001;
mem2[7461] = 10'b0111101001;
mem2[7462] = 10'b0111101001;
mem2[7463] = 10'b0111101001;
mem2[7464] = 10'b0111101001;
mem2[7465] = 10'b0111101001;
mem2[7466] = 10'b0111101001;
mem2[7467] = 10'b0111101001;
mem2[7468] = 10'b0111101001;
mem2[7469] = 10'b0111101001;
mem2[7470] = 10'b0111101010;
mem2[7471] = 10'b0111101010;
mem2[7472] = 10'b0111101010;
mem2[7473] = 10'b0111101010;
mem2[7474] = 10'b0111101010;
mem2[7475] = 10'b0111101010;
mem2[7476] = 10'b0111101010;
mem2[7477] = 10'b0111101010;
mem2[7478] = 10'b0111101010;
mem2[7479] = 10'b0111101011;
mem2[7480] = 10'b0111101011;
mem2[7481] = 10'b0111101011;
mem2[7482] = 10'b0111101011;
mem2[7483] = 10'b0111101011;
mem2[7484] = 10'b0111101011;
mem2[7485] = 10'b0111101011;
mem2[7486] = 10'b0111101011;
mem2[7487] = 10'b0111101011;
mem2[7488] = 10'b0111101011;
mem2[7489] = 10'b0111101100;
mem2[7490] = 10'b0111101100;
mem2[7491] = 10'b0111101100;
mem2[7492] = 10'b0111101100;
mem2[7493] = 10'b0111101100;
mem2[7494] = 10'b0111101100;
mem2[7495] = 10'b0111101100;
mem2[7496] = 10'b0111101100;
mem2[7497] = 10'b0111101100;
mem2[7498] = 10'b0111101100;
mem2[7499] = 10'b0111101101;
mem2[7500] = 10'b0111101101;
mem2[7501] = 10'b0111101101;
mem2[7502] = 10'b0111101101;
mem2[7503] = 10'b0111101101;
mem2[7504] = 10'b0111101101;
mem2[7505] = 10'b0111101101;
mem2[7506] = 10'b0111101101;
mem2[7507] = 10'b0111101101;
mem2[7508] = 10'b0111101110;
mem2[7509] = 10'b0111101110;
mem2[7510] = 10'b0111101110;
mem2[7511] = 10'b0111101110;
mem2[7512] = 10'b0111101110;
mem2[7513] = 10'b0111101110;
mem2[7514] = 10'b0111101110;
mem2[7515] = 10'b0111101110;
mem2[7516] = 10'b0111101110;
mem2[7517] = 10'b0111101110;
mem2[7518] = 10'b0111101111;
mem2[7519] = 10'b0111101111;
mem2[7520] = 10'b0111101111;
mem2[7521] = 10'b0111101111;
mem2[7522] = 10'b0111101111;
mem2[7523] = 10'b0111101111;
mem2[7524] = 10'b0111101111;
mem2[7525] = 10'b0111101111;
mem2[7526] = 10'b0111101111;
mem2[7527] = 10'b0111110000;
mem2[7528] = 10'b0111110000;
mem2[7529] = 10'b0111110000;
mem2[7530] = 10'b0111110000;
mem2[7531] = 10'b0111110000;
mem2[7532] = 10'b0111110000;
mem2[7533] = 10'b0111110000;
mem2[7534] = 10'b0111110000;
mem2[7535] = 10'b0111110000;
mem2[7536] = 10'b0111110000;
mem2[7537] = 10'b0111110001;
mem2[7538] = 10'b0111110001;
mem2[7539] = 10'b0111110001;
mem2[7540] = 10'b0111110001;
mem2[7541] = 10'b0111110001;
mem2[7542] = 10'b0111110001;
mem2[7543] = 10'b0111110001;
mem2[7544] = 10'b0111110001;
mem2[7545] = 10'b0111110001;
mem2[7546] = 10'b0111110010;
mem2[7547] = 10'b0111110010;
mem2[7548] = 10'b0111110010;
mem2[7549] = 10'b0111110010;
mem2[7550] = 10'b0111110010;
mem2[7551] = 10'b0111110010;
mem2[7552] = 10'b0111110010;
mem2[7553] = 10'b0111110010;
mem2[7554] = 10'b0111110010;
mem2[7555] = 10'b0111110010;
mem2[7556] = 10'b0111110011;
mem2[7557] = 10'b0111110011;
mem2[7558] = 10'b0111110011;
mem2[7559] = 10'b0111110011;
mem2[7560] = 10'b0111110011;
mem2[7561] = 10'b0111110011;
mem2[7562] = 10'b0111110011;
mem2[7563] = 10'b0111110011;
mem2[7564] = 10'b0111110011;
mem2[7565] = 10'b0111110100;
mem2[7566] = 10'b0111110100;
mem2[7567] = 10'b0111110100;
mem2[7568] = 10'b0111110100;
mem2[7569] = 10'b0111110100;
mem2[7570] = 10'b0111110100;
mem2[7571] = 10'b0111110100;
mem2[7572] = 10'b0111110100;
mem2[7573] = 10'b0111110100;
mem2[7574] = 10'b0111110100;
mem2[7575] = 10'b0111110101;
mem2[7576] = 10'b0111110101;
mem2[7577] = 10'b0111110101;
mem2[7578] = 10'b0111110101;
mem2[7579] = 10'b0111110101;
mem2[7580] = 10'b0111110101;
mem2[7581] = 10'b0111110101;
mem2[7582] = 10'b0111110101;
mem2[7583] = 10'b0111110101;
mem2[7584] = 10'b0111110101;
mem2[7585] = 10'b0111110110;
mem2[7586] = 10'b0111110110;
mem2[7587] = 10'b0111110110;
mem2[7588] = 10'b0111110110;
mem2[7589] = 10'b0111110110;
mem2[7590] = 10'b0111110110;
mem2[7591] = 10'b0111110110;
mem2[7592] = 10'b0111110110;
mem2[7593] = 10'b0111110110;
mem2[7594] = 10'b0111110111;
mem2[7595] = 10'b0111110111;
mem2[7596] = 10'b0111110111;
mem2[7597] = 10'b0111110111;
mem2[7598] = 10'b0111110111;
mem2[7599] = 10'b0111110111;
mem2[7600] = 10'b0111110111;
mem2[7601] = 10'b0111110111;
mem2[7602] = 10'b0111110111;
mem2[7603] = 10'b0111110111;
mem2[7604] = 10'b0111111000;
mem2[7605] = 10'b0111111000;
mem2[7606] = 10'b0111111000;
mem2[7607] = 10'b0111111000;
mem2[7608] = 10'b0111111000;
mem2[7609] = 10'b0111111000;
mem2[7610] = 10'b0111111000;
mem2[7611] = 10'b0111111000;
mem2[7612] = 10'b0111111000;
mem2[7613] = 10'b0111111001;
mem2[7614] = 10'b0111111001;
mem2[7615] = 10'b0111111001;
mem2[7616] = 10'b0111111001;
mem2[7617] = 10'b0111111001;
mem2[7618] = 10'b0111111001;
mem2[7619] = 10'b0111111001;
mem2[7620] = 10'b0111111001;
mem2[7621] = 10'b0111111001;
mem2[7622] = 10'b0111111001;
mem2[7623] = 10'b0111111010;
mem2[7624] = 10'b0111111010;
mem2[7625] = 10'b0111111010;
mem2[7626] = 10'b0111111010;
mem2[7627] = 10'b0111111010;
mem2[7628] = 10'b0111111010;
mem2[7629] = 10'b0111111010;
mem2[7630] = 10'b0111111010;
mem2[7631] = 10'b0111111010;
mem2[7632] = 10'b0111111011;
mem2[7633] = 10'b0111111011;
mem2[7634] = 10'b0111111011;
mem2[7635] = 10'b0111111011;
mem2[7636] = 10'b0111111011;
mem2[7637] = 10'b0111111011;
mem2[7638] = 10'b0111111011;
mem2[7639] = 10'b0111111011;
mem2[7640] = 10'b0111111011;
mem2[7641] = 10'b0111111011;
mem2[7642] = 10'b0111111100;
mem2[7643] = 10'b0111111100;
mem2[7644] = 10'b0111111100;
mem2[7645] = 10'b0111111100;
mem2[7646] = 10'b0111111100;
mem2[7647] = 10'b0111111100;
mem2[7648] = 10'b0111111100;
mem2[7649] = 10'b0111111100;
mem2[7650] = 10'b0111111100;
mem2[7651] = 10'b0111111101;
mem2[7652] = 10'b0111111101;
mem2[7653] = 10'b0111111101;
mem2[7654] = 10'b0111111101;
mem2[7655] = 10'b0111111101;
mem2[7656] = 10'b0111111101;
mem2[7657] = 10'b0111111101;
mem2[7658] = 10'b0111111101;
mem2[7659] = 10'b0111111101;
mem2[7660] = 10'b0111111101;
mem2[7661] = 10'b0111111110;
mem2[7662] = 10'b0111111110;
mem2[7663] = 10'b0111111110;
mem2[7664] = 10'b0111111110;
mem2[7665] = 10'b0111111110;
mem2[7666] = 10'b0111111110;
mem2[7667] = 10'b0111111110;
mem2[7668] = 10'b0111111110;
mem2[7669] = 10'b0111111110;
mem2[7670] = 10'b0111111111;
mem2[7671] = 10'b0111111111;
mem2[7672] = 10'b0111111111;
mem2[7673] = 10'b0111111111;
mem2[7674] = 10'b0111111111;
mem2[7675] = 10'b0111111111;
mem2[7676] = 10'b0111111111;
mem2[7677] = 10'b0111111111;
mem2[7678] = 10'b0111111111;
mem2[7679] = 10'b0111111111;
mem2[7680] = 10'b1000000000;
mem2[7681] = 10'b1000000000;
mem2[7682] = 10'b1000000000;
mem2[7683] = 10'b1000000000;
mem2[7684] = 10'b1000000000;
mem2[7685] = 10'b1000000000;
mem2[7686] = 10'b1000000000;
mem2[7687] = 10'b1000000000;
mem2[7688] = 10'b1000000000;
mem2[7689] = 10'b1000000000;
mem2[7690] = 10'b1000000001;
mem2[7691] = 10'b1000000001;
mem2[7692] = 10'b1000000001;
mem2[7693] = 10'b1000000001;
mem2[7694] = 10'b1000000001;
mem2[7695] = 10'b1000000001;
mem2[7696] = 10'b1000000001;
mem2[7697] = 10'b1000000001;
mem2[7698] = 10'b1000000001;
mem2[7699] = 10'b1000000010;
mem2[7700] = 10'b1000000010;
mem2[7701] = 10'b1000000010;
mem2[7702] = 10'b1000000010;
mem2[7703] = 10'b1000000010;
mem2[7704] = 10'b1000000010;
mem2[7705] = 10'b1000000010;
mem2[7706] = 10'b1000000010;
mem2[7707] = 10'b1000000010;
mem2[7708] = 10'b1000000010;
mem2[7709] = 10'b1000000011;
mem2[7710] = 10'b1000000011;
mem2[7711] = 10'b1000000011;
mem2[7712] = 10'b1000000011;
mem2[7713] = 10'b1000000011;
mem2[7714] = 10'b1000000011;
mem2[7715] = 10'b1000000011;
mem2[7716] = 10'b1000000011;
mem2[7717] = 10'b1000000011;
mem2[7718] = 10'b1000000100;
mem2[7719] = 10'b1000000100;
mem2[7720] = 10'b1000000100;
mem2[7721] = 10'b1000000100;
mem2[7722] = 10'b1000000100;
mem2[7723] = 10'b1000000100;
mem2[7724] = 10'b1000000100;
mem2[7725] = 10'b1000000100;
mem2[7726] = 10'b1000000100;
mem2[7727] = 10'b1000000100;
mem2[7728] = 10'b1000000101;
mem2[7729] = 10'b1000000101;
mem2[7730] = 10'b1000000101;
mem2[7731] = 10'b1000000101;
mem2[7732] = 10'b1000000101;
mem2[7733] = 10'b1000000101;
mem2[7734] = 10'b1000000101;
mem2[7735] = 10'b1000000101;
mem2[7736] = 10'b1000000101;
mem2[7737] = 10'b1000000110;
mem2[7738] = 10'b1000000110;
mem2[7739] = 10'b1000000110;
mem2[7740] = 10'b1000000110;
mem2[7741] = 10'b1000000110;
mem2[7742] = 10'b1000000110;
mem2[7743] = 10'b1000000110;
mem2[7744] = 10'b1000000110;
mem2[7745] = 10'b1000000110;
mem2[7746] = 10'b1000000110;
mem2[7747] = 10'b1000000111;
mem2[7748] = 10'b1000000111;
mem2[7749] = 10'b1000000111;
mem2[7750] = 10'b1000000111;
mem2[7751] = 10'b1000000111;
mem2[7752] = 10'b1000000111;
mem2[7753] = 10'b1000000111;
mem2[7754] = 10'b1000000111;
mem2[7755] = 10'b1000000111;
mem2[7756] = 10'b1000001000;
mem2[7757] = 10'b1000001000;
mem2[7758] = 10'b1000001000;
mem2[7759] = 10'b1000001000;
mem2[7760] = 10'b1000001000;
mem2[7761] = 10'b1000001000;
mem2[7762] = 10'b1000001000;
mem2[7763] = 10'b1000001000;
mem2[7764] = 10'b1000001000;
mem2[7765] = 10'b1000001000;
mem2[7766] = 10'b1000001001;
mem2[7767] = 10'b1000001001;
mem2[7768] = 10'b1000001001;
mem2[7769] = 10'b1000001001;
mem2[7770] = 10'b1000001001;
mem2[7771] = 10'b1000001001;
mem2[7772] = 10'b1000001001;
mem2[7773] = 10'b1000001001;
mem2[7774] = 10'b1000001001;
mem2[7775] = 10'b1000001010;
mem2[7776] = 10'b1000001010;
mem2[7777] = 10'b1000001010;
mem2[7778] = 10'b1000001010;
mem2[7779] = 10'b1000001010;
mem2[7780] = 10'b1000001010;
mem2[7781] = 10'b1000001010;
mem2[7782] = 10'b1000001010;
mem2[7783] = 10'b1000001010;
mem2[7784] = 10'b1000001010;
mem2[7785] = 10'b1000001011;
mem2[7786] = 10'b1000001011;
mem2[7787] = 10'b1000001011;
mem2[7788] = 10'b1000001011;
mem2[7789] = 10'b1000001011;
mem2[7790] = 10'b1000001011;
mem2[7791] = 10'b1000001011;
mem2[7792] = 10'b1000001011;
mem2[7793] = 10'b1000001011;
mem2[7794] = 10'b1000001011;
mem2[7795] = 10'b1000001100;
mem2[7796] = 10'b1000001100;
mem2[7797] = 10'b1000001100;
mem2[7798] = 10'b1000001100;
mem2[7799] = 10'b1000001100;
mem2[7800] = 10'b1000001100;
mem2[7801] = 10'b1000001100;
mem2[7802] = 10'b1000001100;
mem2[7803] = 10'b1000001100;
mem2[7804] = 10'b1000001101;
mem2[7805] = 10'b1000001101;
mem2[7806] = 10'b1000001101;
mem2[7807] = 10'b1000001101;
mem2[7808] = 10'b1000001101;
mem2[7809] = 10'b1000001101;
mem2[7810] = 10'b1000001101;
mem2[7811] = 10'b1000001101;
mem2[7812] = 10'b1000001101;
mem2[7813] = 10'b1000001101;
mem2[7814] = 10'b1000001110;
mem2[7815] = 10'b1000001110;
mem2[7816] = 10'b1000001110;
mem2[7817] = 10'b1000001110;
mem2[7818] = 10'b1000001110;
mem2[7819] = 10'b1000001110;
mem2[7820] = 10'b1000001110;
mem2[7821] = 10'b1000001110;
mem2[7822] = 10'b1000001110;
mem2[7823] = 10'b1000001111;
mem2[7824] = 10'b1000001111;
mem2[7825] = 10'b1000001111;
mem2[7826] = 10'b1000001111;
mem2[7827] = 10'b1000001111;
mem2[7828] = 10'b1000001111;
mem2[7829] = 10'b1000001111;
mem2[7830] = 10'b1000001111;
mem2[7831] = 10'b1000001111;
mem2[7832] = 10'b1000001111;
mem2[7833] = 10'b1000010000;
mem2[7834] = 10'b1000010000;
mem2[7835] = 10'b1000010000;
mem2[7836] = 10'b1000010000;
mem2[7837] = 10'b1000010000;
mem2[7838] = 10'b1000010000;
mem2[7839] = 10'b1000010000;
mem2[7840] = 10'b1000010000;
mem2[7841] = 10'b1000010000;
mem2[7842] = 10'b1000010001;
mem2[7843] = 10'b1000010001;
mem2[7844] = 10'b1000010001;
mem2[7845] = 10'b1000010001;
mem2[7846] = 10'b1000010001;
mem2[7847] = 10'b1000010001;
mem2[7848] = 10'b1000010001;
mem2[7849] = 10'b1000010001;
mem2[7850] = 10'b1000010001;
mem2[7851] = 10'b1000010001;
mem2[7852] = 10'b1000010010;
mem2[7853] = 10'b1000010010;
mem2[7854] = 10'b1000010010;
mem2[7855] = 10'b1000010010;
mem2[7856] = 10'b1000010010;
mem2[7857] = 10'b1000010010;
mem2[7858] = 10'b1000010010;
mem2[7859] = 10'b1000010010;
mem2[7860] = 10'b1000010010;
mem2[7861] = 10'b1000010011;
mem2[7862] = 10'b1000010011;
mem2[7863] = 10'b1000010011;
mem2[7864] = 10'b1000010011;
mem2[7865] = 10'b1000010011;
mem2[7866] = 10'b1000010011;
mem2[7867] = 10'b1000010011;
mem2[7868] = 10'b1000010011;
mem2[7869] = 10'b1000010011;
mem2[7870] = 10'b1000010011;
mem2[7871] = 10'b1000010100;
mem2[7872] = 10'b1000010100;
mem2[7873] = 10'b1000010100;
mem2[7874] = 10'b1000010100;
mem2[7875] = 10'b1000010100;
mem2[7876] = 10'b1000010100;
mem2[7877] = 10'b1000010100;
mem2[7878] = 10'b1000010100;
mem2[7879] = 10'b1000010100;
mem2[7880] = 10'b1000010100;
mem2[7881] = 10'b1000010101;
mem2[7882] = 10'b1000010101;
mem2[7883] = 10'b1000010101;
mem2[7884] = 10'b1000010101;
mem2[7885] = 10'b1000010101;
mem2[7886] = 10'b1000010101;
mem2[7887] = 10'b1000010101;
mem2[7888] = 10'b1000010101;
mem2[7889] = 10'b1000010101;
mem2[7890] = 10'b1000010110;
mem2[7891] = 10'b1000010110;
mem2[7892] = 10'b1000010110;
mem2[7893] = 10'b1000010110;
mem2[7894] = 10'b1000010110;
mem2[7895] = 10'b1000010110;
mem2[7896] = 10'b1000010110;
mem2[7897] = 10'b1000010110;
mem2[7898] = 10'b1000010110;
mem2[7899] = 10'b1000010110;
mem2[7900] = 10'b1000010111;
mem2[7901] = 10'b1000010111;
mem2[7902] = 10'b1000010111;
mem2[7903] = 10'b1000010111;
mem2[7904] = 10'b1000010111;
mem2[7905] = 10'b1000010111;
mem2[7906] = 10'b1000010111;
mem2[7907] = 10'b1000010111;
mem2[7908] = 10'b1000010111;
mem2[7909] = 10'b1000011000;
mem2[7910] = 10'b1000011000;
mem2[7911] = 10'b1000011000;
mem2[7912] = 10'b1000011000;
mem2[7913] = 10'b1000011000;
mem2[7914] = 10'b1000011000;
mem2[7915] = 10'b1000011000;
mem2[7916] = 10'b1000011000;
mem2[7917] = 10'b1000011000;
mem2[7918] = 10'b1000011000;
mem2[7919] = 10'b1000011001;
mem2[7920] = 10'b1000011001;
mem2[7921] = 10'b1000011001;
mem2[7922] = 10'b1000011001;
mem2[7923] = 10'b1000011001;
mem2[7924] = 10'b1000011001;
mem2[7925] = 10'b1000011001;
mem2[7926] = 10'b1000011001;
mem2[7927] = 10'b1000011001;
mem2[7928] = 10'b1000011010;
mem2[7929] = 10'b1000011010;
mem2[7930] = 10'b1000011010;
mem2[7931] = 10'b1000011010;
mem2[7932] = 10'b1000011010;
mem2[7933] = 10'b1000011010;
mem2[7934] = 10'b1000011010;
mem2[7935] = 10'b1000011010;
mem2[7936] = 10'b1000011010;
mem2[7937] = 10'b1000011010;
mem2[7938] = 10'b1000011011;
mem2[7939] = 10'b1000011011;
mem2[7940] = 10'b1000011011;
mem2[7941] = 10'b1000011011;
mem2[7942] = 10'b1000011011;
mem2[7943] = 10'b1000011011;
mem2[7944] = 10'b1000011011;
mem2[7945] = 10'b1000011011;
mem2[7946] = 10'b1000011011;
mem2[7947] = 10'b1000011011;
mem2[7948] = 10'b1000011100;
mem2[7949] = 10'b1000011100;
mem2[7950] = 10'b1000011100;
mem2[7951] = 10'b1000011100;
mem2[7952] = 10'b1000011100;
mem2[7953] = 10'b1000011100;
mem2[7954] = 10'b1000011100;
mem2[7955] = 10'b1000011100;
mem2[7956] = 10'b1000011100;
mem2[7957] = 10'b1000011101;
mem2[7958] = 10'b1000011101;
mem2[7959] = 10'b1000011101;
mem2[7960] = 10'b1000011101;
mem2[7961] = 10'b1000011101;
mem2[7962] = 10'b1000011101;
mem2[7963] = 10'b1000011101;
mem2[7964] = 10'b1000011101;
mem2[7965] = 10'b1000011101;
mem2[7966] = 10'b1000011101;
mem2[7967] = 10'b1000011110;
mem2[7968] = 10'b1000011110;
mem2[7969] = 10'b1000011110;
mem2[7970] = 10'b1000011110;
mem2[7971] = 10'b1000011110;
mem2[7972] = 10'b1000011110;
mem2[7973] = 10'b1000011110;
mem2[7974] = 10'b1000011110;
mem2[7975] = 10'b1000011110;
mem2[7976] = 10'b1000011111;
mem2[7977] = 10'b1000011111;
mem2[7978] = 10'b1000011111;
mem2[7979] = 10'b1000011111;
mem2[7980] = 10'b1000011111;
mem2[7981] = 10'b1000011111;
mem2[7982] = 10'b1000011111;
mem2[7983] = 10'b1000011111;
mem2[7984] = 10'b1000011111;
mem2[7985] = 10'b1000011111;
mem2[7986] = 10'b1000100000;
mem2[7987] = 10'b1000100000;
mem2[7988] = 10'b1000100000;
mem2[7989] = 10'b1000100000;
mem2[7990] = 10'b1000100000;
mem2[7991] = 10'b1000100000;
mem2[7992] = 10'b1000100000;
mem2[7993] = 10'b1000100000;
mem2[7994] = 10'b1000100000;
mem2[7995] = 10'b1000100001;
mem2[7996] = 10'b1000100001;
mem2[7997] = 10'b1000100001;
mem2[7998] = 10'b1000100001;
mem2[7999] = 10'b1000100001;
mem2[8000] = 10'b1000100001;
mem2[8001] = 10'b1000100001;
mem2[8002] = 10'b1000100001;
mem2[8003] = 10'b1000100001;
mem2[8004] = 10'b1000100001;
mem2[8005] = 10'b1000100010;
mem2[8006] = 10'b1000100010;
mem2[8007] = 10'b1000100010;
mem2[8008] = 10'b1000100010;
mem2[8009] = 10'b1000100010;
mem2[8010] = 10'b1000100010;
mem2[8011] = 10'b1000100010;
mem2[8012] = 10'b1000100010;
mem2[8013] = 10'b1000100010;
mem2[8014] = 10'b1000100011;
mem2[8015] = 10'b1000100011;
mem2[8016] = 10'b1000100011;
mem2[8017] = 10'b1000100011;
mem2[8018] = 10'b1000100011;
mem2[8019] = 10'b1000100011;
mem2[8020] = 10'b1000100011;
mem2[8021] = 10'b1000100011;
mem2[8022] = 10'b1000100011;
mem2[8023] = 10'b1000100011;
mem2[8024] = 10'b1000100100;
mem2[8025] = 10'b1000100100;
mem2[8026] = 10'b1000100100;
mem2[8027] = 10'b1000100100;
mem2[8028] = 10'b1000100100;
mem2[8029] = 10'b1000100100;
mem2[8030] = 10'b1000100100;
mem2[8031] = 10'b1000100100;
mem2[8032] = 10'b1000100100;
mem2[8033] = 10'b1000100100;
mem2[8034] = 10'b1000100101;
mem2[8035] = 10'b1000100101;
mem2[8036] = 10'b1000100101;
mem2[8037] = 10'b1000100101;
mem2[8038] = 10'b1000100101;
mem2[8039] = 10'b1000100101;
mem2[8040] = 10'b1000100101;
mem2[8041] = 10'b1000100101;
mem2[8042] = 10'b1000100101;
mem2[8043] = 10'b1000100110;
mem2[8044] = 10'b1000100110;
mem2[8045] = 10'b1000100110;
mem2[8046] = 10'b1000100110;
mem2[8047] = 10'b1000100110;
mem2[8048] = 10'b1000100110;
mem2[8049] = 10'b1000100110;
mem2[8050] = 10'b1000100110;
mem2[8051] = 10'b1000100110;
mem2[8052] = 10'b1000100110;
mem2[8053] = 10'b1000100111;
mem2[8054] = 10'b1000100111;
mem2[8055] = 10'b1000100111;
mem2[8056] = 10'b1000100111;
mem2[8057] = 10'b1000100111;
mem2[8058] = 10'b1000100111;
mem2[8059] = 10'b1000100111;
mem2[8060] = 10'b1000100111;
mem2[8061] = 10'b1000100111;
mem2[8062] = 10'b1000101000;
mem2[8063] = 10'b1000101000;
mem2[8064] = 10'b1000101000;
mem2[8065] = 10'b1000101000;
mem2[8066] = 10'b1000101000;
mem2[8067] = 10'b1000101000;
mem2[8068] = 10'b1000101000;
mem2[8069] = 10'b1000101000;
mem2[8070] = 10'b1000101000;
mem2[8071] = 10'b1000101000;
mem2[8072] = 10'b1000101001;
mem2[8073] = 10'b1000101001;
mem2[8074] = 10'b1000101001;
mem2[8075] = 10'b1000101001;
mem2[8076] = 10'b1000101001;
mem2[8077] = 10'b1000101001;
mem2[8078] = 10'b1000101001;
mem2[8079] = 10'b1000101001;
mem2[8080] = 10'b1000101001;
mem2[8081] = 10'b1000101001;
mem2[8082] = 10'b1000101010;
mem2[8083] = 10'b1000101010;
mem2[8084] = 10'b1000101010;
mem2[8085] = 10'b1000101010;
mem2[8086] = 10'b1000101010;
mem2[8087] = 10'b1000101010;
mem2[8088] = 10'b1000101010;
mem2[8089] = 10'b1000101010;
mem2[8090] = 10'b1000101010;
mem2[8091] = 10'b1000101011;
mem2[8092] = 10'b1000101011;
mem2[8093] = 10'b1000101011;
mem2[8094] = 10'b1000101011;
mem2[8095] = 10'b1000101011;
mem2[8096] = 10'b1000101011;
mem2[8097] = 10'b1000101011;
mem2[8098] = 10'b1000101011;
mem2[8099] = 10'b1000101011;
mem2[8100] = 10'b1000101011;
mem2[8101] = 10'b1000101100;
mem2[8102] = 10'b1000101100;
mem2[8103] = 10'b1000101100;
mem2[8104] = 10'b1000101100;
mem2[8105] = 10'b1000101100;
mem2[8106] = 10'b1000101100;
mem2[8107] = 10'b1000101100;
mem2[8108] = 10'b1000101100;
mem2[8109] = 10'b1000101100;
mem2[8110] = 10'b1000101101;
mem2[8111] = 10'b1000101101;
mem2[8112] = 10'b1000101101;
mem2[8113] = 10'b1000101101;
mem2[8114] = 10'b1000101101;
mem2[8115] = 10'b1000101101;
mem2[8116] = 10'b1000101101;
mem2[8117] = 10'b1000101101;
mem2[8118] = 10'b1000101101;
mem2[8119] = 10'b1000101101;
mem2[8120] = 10'b1000101110;
mem2[8121] = 10'b1000101110;
mem2[8122] = 10'b1000101110;
mem2[8123] = 10'b1000101110;
mem2[8124] = 10'b1000101110;
mem2[8125] = 10'b1000101110;
mem2[8126] = 10'b1000101110;
mem2[8127] = 10'b1000101110;
mem2[8128] = 10'b1000101110;
mem2[8129] = 10'b1000101111;
mem2[8130] = 10'b1000101111;
mem2[8131] = 10'b1000101111;
mem2[8132] = 10'b1000101111;
mem2[8133] = 10'b1000101111;
mem2[8134] = 10'b1000101111;
mem2[8135] = 10'b1000101111;
mem2[8136] = 10'b1000101111;
mem2[8137] = 10'b1000101111;
mem2[8138] = 10'b1000101111;
mem2[8139] = 10'b1000110000;
mem2[8140] = 10'b1000110000;
mem2[8141] = 10'b1000110000;
mem2[8142] = 10'b1000110000;
mem2[8143] = 10'b1000110000;
mem2[8144] = 10'b1000110000;
mem2[8145] = 10'b1000110000;
mem2[8146] = 10'b1000110000;
mem2[8147] = 10'b1000110000;
mem2[8148] = 10'b1000110000;
mem2[8149] = 10'b1000110001;
mem2[8150] = 10'b1000110001;
mem2[8151] = 10'b1000110001;
mem2[8152] = 10'b1000110001;
mem2[8153] = 10'b1000110001;
mem2[8154] = 10'b1000110001;
mem2[8155] = 10'b1000110001;
mem2[8156] = 10'b1000110001;
mem2[8157] = 10'b1000110001;
mem2[8158] = 10'b1000110010;
mem2[8159] = 10'b1000110010;
mem2[8160] = 10'b1000110010;
mem2[8161] = 10'b1000110010;
mem2[8162] = 10'b1000110010;
mem2[8163] = 10'b1000110010;
mem2[8164] = 10'b1000110010;
mem2[8165] = 10'b1000110010;
mem2[8166] = 10'b1000110010;
mem2[8167] = 10'b1000110010;
mem2[8168] = 10'b1000110011;
mem2[8169] = 10'b1000110011;
mem2[8170] = 10'b1000110011;
mem2[8171] = 10'b1000110011;
mem2[8172] = 10'b1000110011;
mem2[8173] = 10'b1000110011;
mem2[8174] = 10'b1000110011;
mem2[8175] = 10'b1000110011;
mem2[8176] = 10'b1000110011;
mem2[8177] = 10'b1000110100;
mem2[8178] = 10'b1000110100;
mem2[8179] = 10'b1000110100;
mem2[8180] = 10'b1000110100;
mem2[8181] = 10'b1000110100;
mem2[8182] = 10'b1000110100;
mem2[8183] = 10'b1000110100;
mem2[8184] = 10'b1000110100;
mem2[8185] = 10'b1000110100;
mem2[8186] = 10'b1000110100;
mem2[8187] = 10'b1000110101;
mem2[8188] = 10'b1000110101;
mem2[8189] = 10'b1000110101;
mem2[8190] = 10'b1000110101;
mem2[8191] = 10'b1000110101;
mem2[8192] = 10'b1000110101;
mem2[8193] = 10'b1000110101;
mem2[8194] = 10'b1000110101;
mem2[8195] = 10'b1000110101;
mem2[8196] = 10'b1000110101;
mem2[8197] = 10'b1000110110;
mem2[8198] = 10'b1000110110;
mem2[8199] = 10'b1000110110;
mem2[8200] = 10'b1000110110;
mem2[8201] = 10'b1000110110;
mem2[8202] = 10'b1000110110;
mem2[8203] = 10'b1000110110;
mem2[8204] = 10'b1000110110;
mem2[8205] = 10'b1000110110;
mem2[8206] = 10'b1000110111;
mem2[8207] = 10'b1000110111;
mem2[8208] = 10'b1000110111;
mem2[8209] = 10'b1000110111;
mem2[8210] = 10'b1000110111;
mem2[8211] = 10'b1000110111;
mem2[8212] = 10'b1000110111;
mem2[8213] = 10'b1000110111;
mem2[8214] = 10'b1000110111;
mem2[8215] = 10'b1000110111;
mem2[8216] = 10'b1000111000;
mem2[8217] = 10'b1000111000;
mem2[8218] = 10'b1000111000;
mem2[8219] = 10'b1000111000;
mem2[8220] = 10'b1000111000;
mem2[8221] = 10'b1000111000;
mem2[8222] = 10'b1000111000;
mem2[8223] = 10'b1000111000;
mem2[8224] = 10'b1000111000;
mem2[8225] = 10'b1000111001;
mem2[8226] = 10'b1000111001;
mem2[8227] = 10'b1000111001;
mem2[8228] = 10'b1000111001;
mem2[8229] = 10'b1000111001;
mem2[8230] = 10'b1000111001;
mem2[8231] = 10'b1000111001;
mem2[8232] = 10'b1000111001;
mem2[8233] = 10'b1000111001;
mem2[8234] = 10'b1000111001;
mem2[8235] = 10'b1000111010;
mem2[8236] = 10'b1000111010;
mem2[8237] = 10'b1000111010;
mem2[8238] = 10'b1000111010;
mem2[8239] = 10'b1000111010;
mem2[8240] = 10'b1000111010;
mem2[8241] = 10'b1000111010;
mem2[8242] = 10'b1000111010;
mem2[8243] = 10'b1000111010;
mem2[8244] = 10'b1000111010;
mem2[8245] = 10'b1000111011;
mem2[8246] = 10'b1000111011;
mem2[8247] = 10'b1000111011;
mem2[8248] = 10'b1000111011;
mem2[8249] = 10'b1000111011;
mem2[8250] = 10'b1000111011;
mem2[8251] = 10'b1000111011;
mem2[8252] = 10'b1000111011;
mem2[8253] = 10'b1000111011;
mem2[8254] = 10'b1000111100;
mem2[8255] = 10'b1000111100;
mem2[8256] = 10'b1000111100;
mem2[8257] = 10'b1000111100;
mem2[8258] = 10'b1000111100;
mem2[8259] = 10'b1000111100;
mem2[8260] = 10'b1000111100;
mem2[8261] = 10'b1000111100;
mem2[8262] = 10'b1000111100;
mem2[8263] = 10'b1000111100;
mem2[8264] = 10'b1000111101;
mem2[8265] = 10'b1000111101;
mem2[8266] = 10'b1000111101;
mem2[8267] = 10'b1000111101;
mem2[8268] = 10'b1000111101;
mem2[8269] = 10'b1000111101;
mem2[8270] = 10'b1000111101;
mem2[8271] = 10'b1000111101;
mem2[8272] = 10'b1000111101;
mem2[8273] = 10'b1000111110;
mem2[8274] = 10'b1000111110;
mem2[8275] = 10'b1000111110;
mem2[8276] = 10'b1000111110;
mem2[8277] = 10'b1000111110;
mem2[8278] = 10'b1000111110;
mem2[8279] = 10'b1000111110;
mem2[8280] = 10'b1000111110;
mem2[8281] = 10'b1000111110;
mem2[8282] = 10'b1000111110;
mem2[8283] = 10'b1000111111;
mem2[8284] = 10'b1000111111;
mem2[8285] = 10'b1000111111;
mem2[8286] = 10'b1000111111;
mem2[8287] = 10'b1000111111;
mem2[8288] = 10'b1000111111;
mem2[8289] = 10'b1000111111;
mem2[8290] = 10'b1000111111;
mem2[8291] = 10'b1000111111;
mem2[8292] = 10'b1000111111;
mem2[8293] = 10'b1001000000;
mem2[8294] = 10'b1001000000;
mem2[8295] = 10'b1001000000;
mem2[8296] = 10'b1001000000;
mem2[8297] = 10'b1001000000;
mem2[8298] = 10'b1001000000;
mem2[8299] = 10'b1001000000;
mem2[8300] = 10'b1001000000;
mem2[8301] = 10'b1001000000;
mem2[8302] = 10'b1001000001;
mem2[8303] = 10'b1001000001;
mem2[8304] = 10'b1001000001;
mem2[8305] = 10'b1001000001;
mem2[8306] = 10'b1001000001;
mem2[8307] = 10'b1001000001;
mem2[8308] = 10'b1001000001;
mem2[8309] = 10'b1001000001;
mem2[8310] = 10'b1001000001;
mem2[8311] = 10'b1001000001;
mem2[8312] = 10'b1001000010;
mem2[8313] = 10'b1001000010;
mem2[8314] = 10'b1001000010;
mem2[8315] = 10'b1001000010;
mem2[8316] = 10'b1001000010;
mem2[8317] = 10'b1001000010;
mem2[8318] = 10'b1001000010;
mem2[8319] = 10'b1001000010;
mem2[8320] = 10'b1001000010;
mem2[8321] = 10'b1001000010;
mem2[8322] = 10'b1001000011;
mem2[8323] = 10'b1001000011;
mem2[8324] = 10'b1001000011;
mem2[8325] = 10'b1001000011;
mem2[8326] = 10'b1001000011;
mem2[8327] = 10'b1001000011;
mem2[8328] = 10'b1001000011;
mem2[8329] = 10'b1001000011;
mem2[8330] = 10'b1001000011;
mem2[8331] = 10'b1001000100;
mem2[8332] = 10'b1001000100;
mem2[8333] = 10'b1001000100;
mem2[8334] = 10'b1001000100;
mem2[8335] = 10'b1001000100;
mem2[8336] = 10'b1001000100;
mem2[8337] = 10'b1001000100;
mem2[8338] = 10'b1001000100;
mem2[8339] = 10'b1001000100;
mem2[8340] = 10'b1001000100;
mem2[8341] = 10'b1001000101;
mem2[8342] = 10'b1001000101;
mem2[8343] = 10'b1001000101;
mem2[8344] = 10'b1001000101;
mem2[8345] = 10'b1001000101;
mem2[8346] = 10'b1001000101;
mem2[8347] = 10'b1001000101;
mem2[8348] = 10'b1001000101;
mem2[8349] = 10'b1001000101;
mem2[8350] = 10'b1001000101;
mem2[8351] = 10'b1001000110;
mem2[8352] = 10'b1001000110;
mem2[8353] = 10'b1001000110;
mem2[8354] = 10'b1001000110;
mem2[8355] = 10'b1001000110;
mem2[8356] = 10'b1001000110;
mem2[8357] = 10'b1001000110;
mem2[8358] = 10'b1001000110;
mem2[8359] = 10'b1001000110;
mem2[8360] = 10'b1001000111;
mem2[8361] = 10'b1001000111;
mem2[8362] = 10'b1001000111;
mem2[8363] = 10'b1001000111;
mem2[8364] = 10'b1001000111;
mem2[8365] = 10'b1001000111;
mem2[8366] = 10'b1001000111;
mem2[8367] = 10'b1001000111;
mem2[8368] = 10'b1001000111;
mem2[8369] = 10'b1001000111;
mem2[8370] = 10'b1001001000;
mem2[8371] = 10'b1001001000;
mem2[8372] = 10'b1001001000;
mem2[8373] = 10'b1001001000;
mem2[8374] = 10'b1001001000;
mem2[8375] = 10'b1001001000;
mem2[8376] = 10'b1001001000;
mem2[8377] = 10'b1001001000;
mem2[8378] = 10'b1001001000;
mem2[8379] = 10'b1001001001;
mem2[8380] = 10'b1001001001;
mem2[8381] = 10'b1001001001;
mem2[8382] = 10'b1001001001;
mem2[8383] = 10'b1001001001;
mem2[8384] = 10'b1001001001;
mem2[8385] = 10'b1001001001;
mem2[8386] = 10'b1001001001;
mem2[8387] = 10'b1001001001;
mem2[8388] = 10'b1001001001;
mem2[8389] = 10'b1001001010;
mem2[8390] = 10'b1001001010;
mem2[8391] = 10'b1001001010;
mem2[8392] = 10'b1001001010;
mem2[8393] = 10'b1001001010;
mem2[8394] = 10'b1001001010;
mem2[8395] = 10'b1001001010;
mem2[8396] = 10'b1001001010;
mem2[8397] = 10'b1001001010;
mem2[8398] = 10'b1001001010;
mem2[8399] = 10'b1001001011;
mem2[8400] = 10'b1001001011;
mem2[8401] = 10'b1001001011;
mem2[8402] = 10'b1001001011;
mem2[8403] = 10'b1001001011;
mem2[8404] = 10'b1001001011;
mem2[8405] = 10'b1001001011;
mem2[8406] = 10'b1001001011;
mem2[8407] = 10'b1001001011;
mem2[8408] = 10'b1001001100;
mem2[8409] = 10'b1001001100;
mem2[8410] = 10'b1001001100;
mem2[8411] = 10'b1001001100;
mem2[8412] = 10'b1001001100;
mem2[8413] = 10'b1001001100;
mem2[8414] = 10'b1001001100;
mem2[8415] = 10'b1001001100;
mem2[8416] = 10'b1001001100;
mem2[8417] = 10'b1001001100;
mem2[8418] = 10'b1001001101;
mem2[8419] = 10'b1001001101;
mem2[8420] = 10'b1001001101;
mem2[8421] = 10'b1001001101;
mem2[8422] = 10'b1001001101;
mem2[8423] = 10'b1001001101;
mem2[8424] = 10'b1001001101;
mem2[8425] = 10'b1001001101;
mem2[8426] = 10'b1001001101;
mem2[8427] = 10'b1001001101;
mem2[8428] = 10'b1001001110;
mem2[8429] = 10'b1001001110;
mem2[8430] = 10'b1001001110;
mem2[8431] = 10'b1001001110;
mem2[8432] = 10'b1001001110;
mem2[8433] = 10'b1001001110;
mem2[8434] = 10'b1001001110;
mem2[8435] = 10'b1001001110;
mem2[8436] = 10'b1001001110;
mem2[8437] = 10'b1001001111;
mem2[8438] = 10'b1001001111;
mem2[8439] = 10'b1001001111;
mem2[8440] = 10'b1001001111;
mem2[8441] = 10'b1001001111;
mem2[8442] = 10'b1001001111;
mem2[8443] = 10'b1001001111;
mem2[8444] = 10'b1001001111;
mem2[8445] = 10'b1001001111;
mem2[8446] = 10'b1001001111;
mem2[8447] = 10'b1001010000;
mem2[8448] = 10'b1001010000;
mem2[8449] = 10'b1001010000;
mem2[8450] = 10'b1001010000;
mem2[8451] = 10'b1001010000;
mem2[8452] = 10'b1001010000;
mem2[8453] = 10'b1001010000;
mem2[8454] = 10'b1001010000;
mem2[8455] = 10'b1001010000;
mem2[8456] = 10'b1001010000;
mem2[8457] = 10'b1001010001;
mem2[8458] = 10'b1001010001;
mem2[8459] = 10'b1001010001;
mem2[8460] = 10'b1001010001;
mem2[8461] = 10'b1001010001;
mem2[8462] = 10'b1001010001;
mem2[8463] = 10'b1001010001;
mem2[8464] = 10'b1001010001;
mem2[8465] = 10'b1001010001;
mem2[8466] = 10'b1001010010;
mem2[8467] = 10'b1001010010;
mem2[8468] = 10'b1001010010;
mem2[8469] = 10'b1001010010;
mem2[8470] = 10'b1001010010;
mem2[8471] = 10'b1001010010;
mem2[8472] = 10'b1001010010;
mem2[8473] = 10'b1001010010;
mem2[8474] = 10'b1001010010;
mem2[8475] = 10'b1001010010;
mem2[8476] = 10'b1001010011;
mem2[8477] = 10'b1001010011;
mem2[8478] = 10'b1001010011;
mem2[8479] = 10'b1001010011;
mem2[8480] = 10'b1001010011;
mem2[8481] = 10'b1001010011;
mem2[8482] = 10'b1001010011;
mem2[8483] = 10'b1001010011;
mem2[8484] = 10'b1001010011;
mem2[8485] = 10'b1001010011;
mem2[8486] = 10'b1001010100;
mem2[8487] = 10'b1001010100;
mem2[8488] = 10'b1001010100;
mem2[8489] = 10'b1001010100;
mem2[8490] = 10'b1001010100;
mem2[8491] = 10'b1001010100;
mem2[8492] = 10'b1001010100;
mem2[8493] = 10'b1001010100;
mem2[8494] = 10'b1001010100;
mem2[8495] = 10'b1001010101;
mem2[8496] = 10'b1001010101;
mem2[8497] = 10'b1001010101;
mem2[8498] = 10'b1001010101;
mem2[8499] = 10'b1001010101;
mem2[8500] = 10'b1001010101;
mem2[8501] = 10'b1001010101;
mem2[8502] = 10'b1001010101;
mem2[8503] = 10'b1001010101;
mem2[8504] = 10'b1001010101;
mem2[8505] = 10'b1001010110;
mem2[8506] = 10'b1001010110;
mem2[8507] = 10'b1001010110;
mem2[8508] = 10'b1001010110;
mem2[8509] = 10'b1001010110;
mem2[8510] = 10'b1001010110;
mem2[8511] = 10'b1001010110;
mem2[8512] = 10'b1001010110;
mem2[8513] = 10'b1001010110;
mem2[8514] = 10'b1001010110;
mem2[8515] = 10'b1001010111;
mem2[8516] = 10'b1001010111;
mem2[8517] = 10'b1001010111;
mem2[8518] = 10'b1001010111;
mem2[8519] = 10'b1001010111;
mem2[8520] = 10'b1001010111;
mem2[8521] = 10'b1001010111;
mem2[8522] = 10'b1001010111;
mem2[8523] = 10'b1001010111;
mem2[8524] = 10'b1001010111;
mem2[8525] = 10'b1001011000;
mem2[8526] = 10'b1001011000;
mem2[8527] = 10'b1001011000;
mem2[8528] = 10'b1001011000;
mem2[8529] = 10'b1001011000;
mem2[8530] = 10'b1001011000;
mem2[8531] = 10'b1001011000;
mem2[8532] = 10'b1001011000;
mem2[8533] = 10'b1001011000;
mem2[8534] = 10'b1001011001;
mem2[8535] = 10'b1001011001;
mem2[8536] = 10'b1001011001;
mem2[8537] = 10'b1001011001;
mem2[8538] = 10'b1001011001;
mem2[8539] = 10'b1001011001;
mem2[8540] = 10'b1001011001;
mem2[8541] = 10'b1001011001;
mem2[8542] = 10'b1001011001;
mem2[8543] = 10'b1001011001;
mem2[8544] = 10'b1001011010;
mem2[8545] = 10'b1001011010;
mem2[8546] = 10'b1001011010;
mem2[8547] = 10'b1001011010;
mem2[8548] = 10'b1001011010;
mem2[8549] = 10'b1001011010;
mem2[8550] = 10'b1001011010;
mem2[8551] = 10'b1001011010;
mem2[8552] = 10'b1001011010;
mem2[8553] = 10'b1001011010;
mem2[8554] = 10'b1001011011;
mem2[8555] = 10'b1001011011;
mem2[8556] = 10'b1001011011;
mem2[8557] = 10'b1001011011;
mem2[8558] = 10'b1001011011;
mem2[8559] = 10'b1001011011;
mem2[8560] = 10'b1001011011;
mem2[8561] = 10'b1001011011;
mem2[8562] = 10'b1001011011;
mem2[8563] = 10'b1001011100;
mem2[8564] = 10'b1001011100;
mem2[8565] = 10'b1001011100;
mem2[8566] = 10'b1001011100;
mem2[8567] = 10'b1001011100;
mem2[8568] = 10'b1001011100;
mem2[8569] = 10'b1001011100;
mem2[8570] = 10'b1001011100;
mem2[8571] = 10'b1001011100;
mem2[8572] = 10'b1001011100;
mem2[8573] = 10'b1001011101;
mem2[8574] = 10'b1001011101;
mem2[8575] = 10'b1001011101;
mem2[8576] = 10'b1001011101;
mem2[8577] = 10'b1001011101;
mem2[8578] = 10'b1001011101;
mem2[8579] = 10'b1001011101;
mem2[8580] = 10'b1001011101;
mem2[8581] = 10'b1001011101;
mem2[8582] = 10'b1001011101;
mem2[8583] = 10'b1001011110;
mem2[8584] = 10'b1001011110;
mem2[8585] = 10'b1001011110;
mem2[8586] = 10'b1001011110;
mem2[8587] = 10'b1001011110;
mem2[8588] = 10'b1001011110;
mem2[8589] = 10'b1001011110;
mem2[8590] = 10'b1001011110;
mem2[8591] = 10'b1001011110;
mem2[8592] = 10'b1001011111;
mem2[8593] = 10'b1001011111;
mem2[8594] = 10'b1001011111;
mem2[8595] = 10'b1001011111;
mem2[8596] = 10'b1001011111;
mem2[8597] = 10'b1001011111;
mem2[8598] = 10'b1001011111;
mem2[8599] = 10'b1001011111;
mem2[8600] = 10'b1001011111;
mem2[8601] = 10'b1001011111;
mem2[8602] = 10'b1001100000;
mem2[8603] = 10'b1001100000;
mem2[8604] = 10'b1001100000;
mem2[8605] = 10'b1001100000;
mem2[8606] = 10'b1001100000;
mem2[8607] = 10'b1001100000;
mem2[8608] = 10'b1001100000;
mem2[8609] = 10'b1001100000;
mem2[8610] = 10'b1001100000;
mem2[8611] = 10'b1001100000;
mem2[8612] = 10'b1001100001;
mem2[8613] = 10'b1001100001;
mem2[8614] = 10'b1001100001;
mem2[8615] = 10'b1001100001;
mem2[8616] = 10'b1001100001;
mem2[8617] = 10'b1001100001;
mem2[8618] = 10'b1001100001;
mem2[8619] = 10'b1001100001;
mem2[8620] = 10'b1001100001;
mem2[8621] = 10'b1001100001;
mem2[8622] = 10'b1001100010;
mem2[8623] = 10'b1001100010;
mem2[8624] = 10'b1001100010;
mem2[8625] = 10'b1001100010;
mem2[8626] = 10'b1001100010;
mem2[8627] = 10'b1001100010;
mem2[8628] = 10'b1001100010;
mem2[8629] = 10'b1001100010;
mem2[8630] = 10'b1001100010;
mem2[8631] = 10'b1001100011;
mem2[8632] = 10'b1001100011;
mem2[8633] = 10'b1001100011;
mem2[8634] = 10'b1001100011;
mem2[8635] = 10'b1001100011;
mem2[8636] = 10'b1001100011;
mem2[8637] = 10'b1001100011;
mem2[8638] = 10'b1001100011;
mem2[8639] = 10'b1001100011;
mem2[8640] = 10'b1001100011;
mem2[8641] = 10'b1001100100;
mem2[8642] = 10'b1001100100;
mem2[8643] = 10'b1001100100;
mem2[8644] = 10'b1001100100;
mem2[8645] = 10'b1001100100;
mem2[8646] = 10'b1001100100;
mem2[8647] = 10'b1001100100;
mem2[8648] = 10'b1001100100;
mem2[8649] = 10'b1001100100;
mem2[8650] = 10'b1001100100;
mem2[8651] = 10'b1001100101;
mem2[8652] = 10'b1001100101;
mem2[8653] = 10'b1001100101;
mem2[8654] = 10'b1001100101;
mem2[8655] = 10'b1001100101;
mem2[8656] = 10'b1001100101;
mem2[8657] = 10'b1001100101;
mem2[8658] = 10'b1001100101;
mem2[8659] = 10'b1001100101;
mem2[8660] = 10'b1001100101;
mem2[8661] = 10'b1001100110;
mem2[8662] = 10'b1001100110;
mem2[8663] = 10'b1001100110;
mem2[8664] = 10'b1001100110;
mem2[8665] = 10'b1001100110;
mem2[8666] = 10'b1001100110;
mem2[8667] = 10'b1001100110;
mem2[8668] = 10'b1001100110;
mem2[8669] = 10'b1001100110;
mem2[8670] = 10'b1001100111;
mem2[8671] = 10'b1001100111;
mem2[8672] = 10'b1001100111;
mem2[8673] = 10'b1001100111;
mem2[8674] = 10'b1001100111;
mem2[8675] = 10'b1001100111;
mem2[8676] = 10'b1001100111;
mem2[8677] = 10'b1001100111;
mem2[8678] = 10'b1001100111;
mem2[8679] = 10'b1001100111;
mem2[8680] = 10'b1001101000;
mem2[8681] = 10'b1001101000;
mem2[8682] = 10'b1001101000;
mem2[8683] = 10'b1001101000;
mem2[8684] = 10'b1001101000;
mem2[8685] = 10'b1001101000;
mem2[8686] = 10'b1001101000;
mem2[8687] = 10'b1001101000;
mem2[8688] = 10'b1001101000;
mem2[8689] = 10'b1001101000;
mem2[8690] = 10'b1001101001;
mem2[8691] = 10'b1001101001;
mem2[8692] = 10'b1001101001;
mem2[8693] = 10'b1001101001;
mem2[8694] = 10'b1001101001;
mem2[8695] = 10'b1001101001;
mem2[8696] = 10'b1001101001;
mem2[8697] = 10'b1001101001;
mem2[8698] = 10'b1001101001;
mem2[8699] = 10'b1001101001;
mem2[8700] = 10'b1001101010;
mem2[8701] = 10'b1001101010;
mem2[8702] = 10'b1001101010;
mem2[8703] = 10'b1001101010;
mem2[8704] = 10'b1001101010;
mem2[8705] = 10'b1001101010;
mem2[8706] = 10'b1001101010;
mem2[8707] = 10'b1001101010;
mem2[8708] = 10'b1001101010;
mem2[8709] = 10'b1001101011;
mem2[8710] = 10'b1001101011;
mem2[8711] = 10'b1001101011;
mem2[8712] = 10'b1001101011;
mem2[8713] = 10'b1001101011;
mem2[8714] = 10'b1001101011;
mem2[8715] = 10'b1001101011;
mem2[8716] = 10'b1001101011;
mem2[8717] = 10'b1001101011;
mem2[8718] = 10'b1001101011;
mem2[8719] = 10'b1001101100;
mem2[8720] = 10'b1001101100;
mem2[8721] = 10'b1001101100;
mem2[8722] = 10'b1001101100;
mem2[8723] = 10'b1001101100;
mem2[8724] = 10'b1001101100;
mem2[8725] = 10'b1001101100;
mem2[8726] = 10'b1001101100;
mem2[8727] = 10'b1001101100;
mem2[8728] = 10'b1001101100;
mem2[8729] = 10'b1001101101;
mem2[8730] = 10'b1001101101;
mem2[8731] = 10'b1001101101;
mem2[8732] = 10'b1001101101;
mem2[8733] = 10'b1001101101;
mem2[8734] = 10'b1001101101;
mem2[8735] = 10'b1001101101;
mem2[8736] = 10'b1001101101;
mem2[8737] = 10'b1001101101;
mem2[8738] = 10'b1001101101;
mem2[8739] = 10'b1001101110;
mem2[8740] = 10'b1001101110;
mem2[8741] = 10'b1001101110;
mem2[8742] = 10'b1001101110;
mem2[8743] = 10'b1001101110;
mem2[8744] = 10'b1001101110;
mem2[8745] = 10'b1001101110;
mem2[8746] = 10'b1001101110;
mem2[8747] = 10'b1001101110;
mem2[8748] = 10'b1001101111;
mem2[8749] = 10'b1001101111;
mem2[8750] = 10'b1001101111;
mem2[8751] = 10'b1001101111;
mem2[8752] = 10'b1001101111;
mem2[8753] = 10'b1001101111;
mem2[8754] = 10'b1001101111;
mem2[8755] = 10'b1001101111;
mem2[8756] = 10'b1001101111;
mem2[8757] = 10'b1001101111;
mem2[8758] = 10'b1001110000;
mem2[8759] = 10'b1001110000;
mem2[8760] = 10'b1001110000;
mem2[8761] = 10'b1001110000;
mem2[8762] = 10'b1001110000;
mem2[8763] = 10'b1001110000;
mem2[8764] = 10'b1001110000;
mem2[8765] = 10'b1001110000;
mem2[8766] = 10'b1001110000;
mem2[8767] = 10'b1001110000;
mem2[8768] = 10'b1001110001;
mem2[8769] = 10'b1001110001;
mem2[8770] = 10'b1001110001;
mem2[8771] = 10'b1001110001;
mem2[8772] = 10'b1001110001;
mem2[8773] = 10'b1001110001;
mem2[8774] = 10'b1001110001;
mem2[8775] = 10'b1001110001;
mem2[8776] = 10'b1001110001;
mem2[8777] = 10'b1001110001;
mem2[8778] = 10'b1001110010;
mem2[8779] = 10'b1001110010;
mem2[8780] = 10'b1001110010;
mem2[8781] = 10'b1001110010;
mem2[8782] = 10'b1001110010;
mem2[8783] = 10'b1001110010;
mem2[8784] = 10'b1001110010;
mem2[8785] = 10'b1001110010;
mem2[8786] = 10'b1001110010;
mem2[8787] = 10'b1001110010;
mem2[8788] = 10'b1001110011;
mem2[8789] = 10'b1001110011;
mem2[8790] = 10'b1001110011;
mem2[8791] = 10'b1001110011;
mem2[8792] = 10'b1001110011;
mem2[8793] = 10'b1001110011;
mem2[8794] = 10'b1001110011;
mem2[8795] = 10'b1001110011;
mem2[8796] = 10'b1001110011;
mem2[8797] = 10'b1001110100;
mem2[8798] = 10'b1001110100;
mem2[8799] = 10'b1001110100;
mem2[8800] = 10'b1001110100;
mem2[8801] = 10'b1001110100;
mem2[8802] = 10'b1001110100;
mem2[8803] = 10'b1001110100;
mem2[8804] = 10'b1001110100;
mem2[8805] = 10'b1001110100;
mem2[8806] = 10'b1001110100;
mem2[8807] = 10'b1001110101;
mem2[8808] = 10'b1001110101;
mem2[8809] = 10'b1001110101;
mem2[8810] = 10'b1001110101;
mem2[8811] = 10'b1001110101;
mem2[8812] = 10'b1001110101;
mem2[8813] = 10'b1001110101;
mem2[8814] = 10'b1001110101;
mem2[8815] = 10'b1001110101;
mem2[8816] = 10'b1001110101;
mem2[8817] = 10'b1001110110;
mem2[8818] = 10'b1001110110;
mem2[8819] = 10'b1001110110;
mem2[8820] = 10'b1001110110;
mem2[8821] = 10'b1001110110;
mem2[8822] = 10'b1001110110;
mem2[8823] = 10'b1001110110;
mem2[8824] = 10'b1001110110;
mem2[8825] = 10'b1001110110;
mem2[8826] = 10'b1001110110;
mem2[8827] = 10'b1001110111;
mem2[8828] = 10'b1001110111;
mem2[8829] = 10'b1001110111;
mem2[8830] = 10'b1001110111;
mem2[8831] = 10'b1001110111;
mem2[8832] = 10'b1001110111;
mem2[8833] = 10'b1001110111;
mem2[8834] = 10'b1001110111;
mem2[8835] = 10'b1001110111;
mem2[8836] = 10'b1001110111;
mem2[8837] = 10'b1001111000;
mem2[8838] = 10'b1001111000;
mem2[8839] = 10'b1001111000;
mem2[8840] = 10'b1001111000;
mem2[8841] = 10'b1001111000;
mem2[8842] = 10'b1001111000;
mem2[8843] = 10'b1001111000;
mem2[8844] = 10'b1001111000;
mem2[8845] = 10'b1001111000;
mem2[8846] = 10'b1001111001;
mem2[8847] = 10'b1001111001;
mem2[8848] = 10'b1001111001;
mem2[8849] = 10'b1001111001;
mem2[8850] = 10'b1001111001;
mem2[8851] = 10'b1001111001;
mem2[8852] = 10'b1001111001;
mem2[8853] = 10'b1001111001;
mem2[8854] = 10'b1001111001;
mem2[8855] = 10'b1001111001;
mem2[8856] = 10'b1001111010;
mem2[8857] = 10'b1001111010;
mem2[8858] = 10'b1001111010;
mem2[8859] = 10'b1001111010;
mem2[8860] = 10'b1001111010;
mem2[8861] = 10'b1001111010;
mem2[8862] = 10'b1001111010;
mem2[8863] = 10'b1001111010;
mem2[8864] = 10'b1001111010;
mem2[8865] = 10'b1001111010;
mem2[8866] = 10'b1001111011;
mem2[8867] = 10'b1001111011;
mem2[8868] = 10'b1001111011;
mem2[8869] = 10'b1001111011;
mem2[8870] = 10'b1001111011;
mem2[8871] = 10'b1001111011;
mem2[8872] = 10'b1001111011;
mem2[8873] = 10'b1001111011;
mem2[8874] = 10'b1001111011;
mem2[8875] = 10'b1001111011;
mem2[8876] = 10'b1001111100;
mem2[8877] = 10'b1001111100;
mem2[8878] = 10'b1001111100;
mem2[8879] = 10'b1001111100;
mem2[8880] = 10'b1001111100;
mem2[8881] = 10'b1001111100;
mem2[8882] = 10'b1001111100;
mem2[8883] = 10'b1001111100;
mem2[8884] = 10'b1001111100;
mem2[8885] = 10'b1001111100;
mem2[8886] = 10'b1001111101;
mem2[8887] = 10'b1001111101;
mem2[8888] = 10'b1001111101;
mem2[8889] = 10'b1001111101;
mem2[8890] = 10'b1001111101;
mem2[8891] = 10'b1001111101;
mem2[8892] = 10'b1001111101;
mem2[8893] = 10'b1001111101;
mem2[8894] = 10'b1001111101;
mem2[8895] = 10'b1001111101;
mem2[8896] = 10'b1001111110;
mem2[8897] = 10'b1001111110;
mem2[8898] = 10'b1001111110;
mem2[8899] = 10'b1001111110;
mem2[8900] = 10'b1001111110;
mem2[8901] = 10'b1001111110;
mem2[8902] = 10'b1001111110;
mem2[8903] = 10'b1001111110;
mem2[8904] = 10'b1001111110;
mem2[8905] = 10'b1001111110;
mem2[8906] = 10'b1001111111;
mem2[8907] = 10'b1001111111;
mem2[8908] = 10'b1001111111;
mem2[8909] = 10'b1001111111;
mem2[8910] = 10'b1001111111;
mem2[8911] = 10'b1001111111;
mem2[8912] = 10'b1001111111;
mem2[8913] = 10'b1001111111;
mem2[8914] = 10'b1001111111;
mem2[8915] = 10'b1010000000;
mem2[8916] = 10'b1010000000;
mem2[8917] = 10'b1010000000;
mem2[8918] = 10'b1010000000;
mem2[8919] = 10'b1010000000;
mem2[8920] = 10'b1010000000;
mem2[8921] = 10'b1010000000;
mem2[8922] = 10'b1010000000;
mem2[8923] = 10'b1010000000;
mem2[8924] = 10'b1010000000;
mem2[8925] = 10'b1010000001;
mem2[8926] = 10'b1010000001;
mem2[8927] = 10'b1010000001;
mem2[8928] = 10'b1010000001;
mem2[8929] = 10'b1010000001;
mem2[8930] = 10'b1010000001;
mem2[8931] = 10'b1010000001;
mem2[8932] = 10'b1010000001;
mem2[8933] = 10'b1010000001;
mem2[8934] = 10'b1010000001;
mem2[8935] = 10'b1010000010;
mem2[8936] = 10'b1010000010;
mem2[8937] = 10'b1010000010;
mem2[8938] = 10'b1010000010;
mem2[8939] = 10'b1010000010;
mem2[8940] = 10'b1010000010;
mem2[8941] = 10'b1010000010;
mem2[8942] = 10'b1010000010;
mem2[8943] = 10'b1010000010;
mem2[8944] = 10'b1010000010;
mem2[8945] = 10'b1010000011;
mem2[8946] = 10'b1010000011;
mem2[8947] = 10'b1010000011;
mem2[8948] = 10'b1010000011;
mem2[8949] = 10'b1010000011;
mem2[8950] = 10'b1010000011;
mem2[8951] = 10'b1010000011;
mem2[8952] = 10'b1010000011;
mem2[8953] = 10'b1010000011;
mem2[8954] = 10'b1010000011;
mem2[8955] = 10'b1010000100;
mem2[8956] = 10'b1010000100;
mem2[8957] = 10'b1010000100;
mem2[8958] = 10'b1010000100;
mem2[8959] = 10'b1010000100;
mem2[8960] = 10'b1010000100;
mem2[8961] = 10'b1010000100;
mem2[8962] = 10'b1010000100;
mem2[8963] = 10'b1010000100;
mem2[8964] = 10'b1010000100;
mem2[8965] = 10'b1010000101;
mem2[8966] = 10'b1010000101;
mem2[8967] = 10'b1010000101;
mem2[8968] = 10'b1010000101;
mem2[8969] = 10'b1010000101;
mem2[8970] = 10'b1010000101;
mem2[8971] = 10'b1010000101;
mem2[8972] = 10'b1010000101;
mem2[8973] = 10'b1010000101;
mem2[8974] = 10'b1010000101;
mem2[8975] = 10'b1010000110;
mem2[8976] = 10'b1010000110;
mem2[8977] = 10'b1010000110;
mem2[8978] = 10'b1010000110;
mem2[8979] = 10'b1010000110;
mem2[8980] = 10'b1010000110;
mem2[8981] = 10'b1010000110;
mem2[8982] = 10'b1010000110;
mem2[8983] = 10'b1010000110;
mem2[8984] = 10'b1010000110;
mem2[8985] = 10'b1010000111;
mem2[8986] = 10'b1010000111;
mem2[8987] = 10'b1010000111;
mem2[8988] = 10'b1010000111;
mem2[8989] = 10'b1010000111;
mem2[8990] = 10'b1010000111;
mem2[8991] = 10'b1010000111;
mem2[8992] = 10'b1010000111;
mem2[8993] = 10'b1010000111;
mem2[8994] = 10'b1010001000;
mem2[8995] = 10'b1010001000;
mem2[8996] = 10'b1010001000;
mem2[8997] = 10'b1010001000;
mem2[8998] = 10'b1010001000;
mem2[8999] = 10'b1010001000;
mem2[9000] = 10'b1010001000;
mem2[9001] = 10'b1010001000;
mem2[9002] = 10'b1010001000;
mem2[9003] = 10'b1010001000;
mem2[9004] = 10'b1010001001;
mem2[9005] = 10'b1010001001;
mem2[9006] = 10'b1010001001;
mem2[9007] = 10'b1010001001;
mem2[9008] = 10'b1010001001;
mem2[9009] = 10'b1010001001;
mem2[9010] = 10'b1010001001;
mem2[9011] = 10'b1010001001;
mem2[9012] = 10'b1010001001;
mem2[9013] = 10'b1010001001;
mem2[9014] = 10'b1010001010;
mem2[9015] = 10'b1010001010;
mem2[9016] = 10'b1010001010;
mem2[9017] = 10'b1010001010;
mem2[9018] = 10'b1010001010;
mem2[9019] = 10'b1010001010;
mem2[9020] = 10'b1010001010;
mem2[9021] = 10'b1010001010;
mem2[9022] = 10'b1010001010;
mem2[9023] = 10'b1010001010;
mem2[9024] = 10'b1010001011;
mem2[9025] = 10'b1010001011;
mem2[9026] = 10'b1010001011;
mem2[9027] = 10'b1010001011;
mem2[9028] = 10'b1010001011;
mem2[9029] = 10'b1010001011;
mem2[9030] = 10'b1010001011;
mem2[9031] = 10'b1010001011;
mem2[9032] = 10'b1010001011;
mem2[9033] = 10'b1010001011;
mem2[9034] = 10'b1010001100;
mem2[9035] = 10'b1010001100;
mem2[9036] = 10'b1010001100;
mem2[9037] = 10'b1010001100;
mem2[9038] = 10'b1010001100;
mem2[9039] = 10'b1010001100;
mem2[9040] = 10'b1010001100;
mem2[9041] = 10'b1010001100;
mem2[9042] = 10'b1010001100;
mem2[9043] = 10'b1010001100;
mem2[9044] = 10'b1010001101;
mem2[9045] = 10'b1010001101;
mem2[9046] = 10'b1010001101;
mem2[9047] = 10'b1010001101;
mem2[9048] = 10'b1010001101;
mem2[9049] = 10'b1010001101;
mem2[9050] = 10'b1010001101;
mem2[9051] = 10'b1010001101;
mem2[9052] = 10'b1010001101;
mem2[9053] = 10'b1010001101;
mem2[9054] = 10'b1010001110;
mem2[9055] = 10'b1010001110;
mem2[9056] = 10'b1010001110;
mem2[9057] = 10'b1010001110;
mem2[9058] = 10'b1010001110;
mem2[9059] = 10'b1010001110;
mem2[9060] = 10'b1010001110;
mem2[9061] = 10'b1010001110;
mem2[9062] = 10'b1010001110;
mem2[9063] = 10'b1010001110;
mem2[9064] = 10'b1010001111;
mem2[9065] = 10'b1010001111;
mem2[9066] = 10'b1010001111;
mem2[9067] = 10'b1010001111;
mem2[9068] = 10'b1010001111;
mem2[9069] = 10'b1010001111;
mem2[9070] = 10'b1010001111;
mem2[9071] = 10'b1010001111;
mem2[9072] = 10'b1010001111;
mem2[9073] = 10'b1010001111;
mem2[9074] = 10'b1010010000;
mem2[9075] = 10'b1010010000;
mem2[9076] = 10'b1010010000;
mem2[9077] = 10'b1010010000;
mem2[9078] = 10'b1010010000;
mem2[9079] = 10'b1010010000;
mem2[9080] = 10'b1010010000;
mem2[9081] = 10'b1010010000;
mem2[9082] = 10'b1010010000;
mem2[9083] = 10'b1010010000;
mem2[9084] = 10'b1010010001;
mem2[9085] = 10'b1010010001;
mem2[9086] = 10'b1010010001;
mem2[9087] = 10'b1010010001;
mem2[9088] = 10'b1010010001;
mem2[9089] = 10'b1010010001;
mem2[9090] = 10'b1010010001;
mem2[9091] = 10'b1010010001;
mem2[9092] = 10'b1010010001;
mem2[9093] = 10'b1010010001;
mem2[9094] = 10'b1010010010;
mem2[9095] = 10'b1010010010;
mem2[9096] = 10'b1010010010;
mem2[9097] = 10'b1010010010;
mem2[9098] = 10'b1010010010;
mem2[9099] = 10'b1010010010;
mem2[9100] = 10'b1010010010;
mem2[9101] = 10'b1010010010;
mem2[9102] = 10'b1010010010;
mem2[9103] = 10'b1010010010;
mem2[9104] = 10'b1010010011;
mem2[9105] = 10'b1010010011;
mem2[9106] = 10'b1010010011;
mem2[9107] = 10'b1010010011;
mem2[9108] = 10'b1010010011;
mem2[9109] = 10'b1010010011;
mem2[9110] = 10'b1010010011;
mem2[9111] = 10'b1010010011;
mem2[9112] = 10'b1010010011;
mem2[9113] = 10'b1010010011;
mem2[9114] = 10'b1010010100;
mem2[9115] = 10'b1010010100;
mem2[9116] = 10'b1010010100;
mem2[9117] = 10'b1010010100;
mem2[9118] = 10'b1010010100;
mem2[9119] = 10'b1010010100;
mem2[9120] = 10'b1010010100;
mem2[9121] = 10'b1010010100;
mem2[9122] = 10'b1010010100;
mem2[9123] = 10'b1010010100;
mem2[9124] = 10'b1010010101;
mem2[9125] = 10'b1010010101;
mem2[9126] = 10'b1010010101;
mem2[9127] = 10'b1010010101;
mem2[9128] = 10'b1010010101;
mem2[9129] = 10'b1010010101;
mem2[9130] = 10'b1010010101;
mem2[9131] = 10'b1010010101;
mem2[9132] = 10'b1010010101;
mem2[9133] = 10'b1010010101;
mem2[9134] = 10'b1010010110;
mem2[9135] = 10'b1010010110;
mem2[9136] = 10'b1010010110;
mem2[9137] = 10'b1010010110;
mem2[9138] = 10'b1010010110;
mem2[9139] = 10'b1010010110;
mem2[9140] = 10'b1010010110;
mem2[9141] = 10'b1010010110;
mem2[9142] = 10'b1010010110;
mem2[9143] = 10'b1010010110;
mem2[9144] = 10'b1010010111;
mem2[9145] = 10'b1010010111;
mem2[9146] = 10'b1010010111;
mem2[9147] = 10'b1010010111;
mem2[9148] = 10'b1010010111;
mem2[9149] = 10'b1010010111;
mem2[9150] = 10'b1010010111;
mem2[9151] = 10'b1010010111;
mem2[9152] = 10'b1010010111;
mem2[9153] = 10'b1010010111;
mem2[9154] = 10'b1010011000;
mem2[9155] = 10'b1010011000;
mem2[9156] = 10'b1010011000;
mem2[9157] = 10'b1010011000;
mem2[9158] = 10'b1010011000;
mem2[9159] = 10'b1010011000;
mem2[9160] = 10'b1010011000;
mem2[9161] = 10'b1010011000;
mem2[9162] = 10'b1010011000;
mem2[9163] = 10'b1010011000;
mem2[9164] = 10'b1010011001;
mem2[9165] = 10'b1010011001;
mem2[9166] = 10'b1010011001;
mem2[9167] = 10'b1010011001;
mem2[9168] = 10'b1010011001;
mem2[9169] = 10'b1010011001;
mem2[9170] = 10'b1010011001;
mem2[9171] = 10'b1010011001;
mem2[9172] = 10'b1010011001;
mem2[9173] = 10'b1010011001;
mem2[9174] = 10'b1010011010;
mem2[9175] = 10'b1010011010;
mem2[9176] = 10'b1010011010;
mem2[9177] = 10'b1010011010;
mem2[9178] = 10'b1010011010;
mem2[9179] = 10'b1010011010;
mem2[9180] = 10'b1010011010;
mem2[9181] = 10'b1010011010;
mem2[9182] = 10'b1010011010;
mem2[9183] = 10'b1010011010;
mem2[9184] = 10'b1010011011;
mem2[9185] = 10'b1010011011;
mem2[9186] = 10'b1010011011;
mem2[9187] = 10'b1010011011;
mem2[9188] = 10'b1010011011;
mem2[9189] = 10'b1010011011;
mem2[9190] = 10'b1010011011;
mem2[9191] = 10'b1010011011;
mem2[9192] = 10'b1010011011;
mem2[9193] = 10'b1010011011;
mem2[9194] = 10'b1010011100;
mem2[9195] = 10'b1010011100;
mem2[9196] = 10'b1010011100;
mem2[9197] = 10'b1010011100;
mem2[9198] = 10'b1010011100;
mem2[9199] = 10'b1010011100;
mem2[9200] = 10'b1010011100;
mem2[9201] = 10'b1010011100;
mem2[9202] = 10'b1010011100;
mem2[9203] = 10'b1010011100;
mem2[9204] = 10'b1010011101;
mem2[9205] = 10'b1010011101;
mem2[9206] = 10'b1010011101;
mem2[9207] = 10'b1010011101;
mem2[9208] = 10'b1010011101;
mem2[9209] = 10'b1010011101;
mem2[9210] = 10'b1010011101;
mem2[9211] = 10'b1010011101;
mem2[9212] = 10'b1010011101;
mem2[9213] = 10'b1010011101;
mem2[9214] = 10'b1010011110;
mem2[9215] = 10'b1010011110;
mem2[9216] = 10'b1010011110;
mem2[9217] = 10'b1010011110;
mem2[9218] = 10'b1010011110;
mem2[9219] = 10'b1010011110;
mem2[9220] = 10'b1010011110;
mem2[9221] = 10'b1010011110;
mem2[9222] = 10'b1010011110;
mem2[9223] = 10'b1010011110;
mem2[9224] = 10'b1010011111;
mem2[9225] = 10'b1010011111;
mem2[9226] = 10'b1010011111;
mem2[9227] = 10'b1010011111;
mem2[9228] = 10'b1010011111;
mem2[9229] = 10'b1010011111;
mem2[9230] = 10'b1010011111;
mem2[9231] = 10'b1010011111;
mem2[9232] = 10'b1010011111;
mem2[9233] = 10'b1010011111;
mem2[9234] = 10'b1010100000;
mem2[9235] = 10'b1010100000;
mem2[9236] = 10'b1010100000;
mem2[9237] = 10'b1010100000;
mem2[9238] = 10'b1010100000;
mem2[9239] = 10'b1010100000;
mem2[9240] = 10'b1010100000;
mem2[9241] = 10'b1010100000;
mem2[9242] = 10'b1010100000;
mem2[9243] = 10'b1010100000;
mem2[9244] = 10'b1010100001;
mem2[9245] = 10'b1010100001;
mem2[9246] = 10'b1010100001;
mem2[9247] = 10'b1010100001;
mem2[9248] = 10'b1010100001;
mem2[9249] = 10'b1010100001;
mem2[9250] = 10'b1010100001;
mem2[9251] = 10'b1010100001;
mem2[9252] = 10'b1010100001;
mem2[9253] = 10'b1010100001;
mem2[9254] = 10'b1010100010;
mem2[9255] = 10'b1010100010;
mem2[9256] = 10'b1010100010;
mem2[9257] = 10'b1010100010;
mem2[9258] = 10'b1010100010;
mem2[9259] = 10'b1010100010;
mem2[9260] = 10'b1010100010;
mem2[9261] = 10'b1010100010;
mem2[9262] = 10'b1010100010;
mem2[9263] = 10'b1010100010;
mem2[9264] = 10'b1010100011;
mem2[9265] = 10'b1010100011;
mem2[9266] = 10'b1010100011;
mem2[9267] = 10'b1010100011;
mem2[9268] = 10'b1010100011;
mem2[9269] = 10'b1010100011;
mem2[9270] = 10'b1010100011;
mem2[9271] = 10'b1010100011;
mem2[9272] = 10'b1010100011;
mem2[9273] = 10'b1010100011;
mem2[9274] = 10'b1010100100;
mem2[9275] = 10'b1010100100;
mem2[9276] = 10'b1010100100;
mem2[9277] = 10'b1010100100;
mem2[9278] = 10'b1010100100;
mem2[9279] = 10'b1010100100;
mem2[9280] = 10'b1010100100;
mem2[9281] = 10'b1010100100;
mem2[9282] = 10'b1010100100;
mem2[9283] = 10'b1010100100;
mem2[9284] = 10'b1010100101;
mem2[9285] = 10'b1010100101;
mem2[9286] = 10'b1010100101;
mem2[9287] = 10'b1010100101;
mem2[9288] = 10'b1010100101;
mem2[9289] = 10'b1010100101;
mem2[9290] = 10'b1010100101;
mem2[9291] = 10'b1010100101;
mem2[9292] = 10'b1010100101;
mem2[9293] = 10'b1010100101;
mem2[9294] = 10'b1010100110;
mem2[9295] = 10'b1010100110;
mem2[9296] = 10'b1010100110;
mem2[9297] = 10'b1010100110;
mem2[9298] = 10'b1010100110;
mem2[9299] = 10'b1010100110;
mem2[9300] = 10'b1010100110;
mem2[9301] = 10'b1010100110;
mem2[9302] = 10'b1010100110;
mem2[9303] = 10'b1010100110;
mem2[9304] = 10'b1010100111;
mem2[9305] = 10'b1010100111;
mem2[9306] = 10'b1010100111;
mem2[9307] = 10'b1010100111;
mem2[9308] = 10'b1010100111;
mem2[9309] = 10'b1010100111;
mem2[9310] = 10'b1010100111;
mem2[9311] = 10'b1010100111;
mem2[9312] = 10'b1010100111;
mem2[9313] = 10'b1010100111;
mem2[9314] = 10'b1010100111;
mem2[9315] = 10'b1010101000;
mem2[9316] = 10'b1010101000;
mem2[9317] = 10'b1010101000;
mem2[9318] = 10'b1010101000;
mem2[9319] = 10'b1010101000;
mem2[9320] = 10'b1010101000;
mem2[9321] = 10'b1010101000;
mem2[9322] = 10'b1010101000;
mem2[9323] = 10'b1010101000;
mem2[9324] = 10'b1010101000;
mem2[9325] = 10'b1010101001;
mem2[9326] = 10'b1010101001;
mem2[9327] = 10'b1010101001;
mem2[9328] = 10'b1010101001;
mem2[9329] = 10'b1010101001;
mem2[9330] = 10'b1010101001;
mem2[9331] = 10'b1010101001;
mem2[9332] = 10'b1010101001;
mem2[9333] = 10'b1010101001;
mem2[9334] = 10'b1010101001;
mem2[9335] = 10'b1010101010;
mem2[9336] = 10'b1010101010;
mem2[9337] = 10'b1010101010;
mem2[9338] = 10'b1010101010;
mem2[9339] = 10'b1010101010;
mem2[9340] = 10'b1010101010;
mem2[9341] = 10'b1010101010;
mem2[9342] = 10'b1010101010;
mem2[9343] = 10'b1010101010;
mem2[9344] = 10'b1010101010;
mem2[9345] = 10'b1010101011;
mem2[9346] = 10'b1010101011;
mem2[9347] = 10'b1010101011;
mem2[9348] = 10'b1010101011;
mem2[9349] = 10'b1010101011;
mem2[9350] = 10'b1010101011;
mem2[9351] = 10'b1010101011;
mem2[9352] = 10'b1010101011;
mem2[9353] = 10'b1010101011;
mem2[9354] = 10'b1010101011;
mem2[9355] = 10'b1010101100;
mem2[9356] = 10'b1010101100;
mem2[9357] = 10'b1010101100;
mem2[9358] = 10'b1010101100;
mem2[9359] = 10'b1010101100;
mem2[9360] = 10'b1010101100;
mem2[9361] = 10'b1010101100;
mem2[9362] = 10'b1010101100;
mem2[9363] = 10'b1010101100;
mem2[9364] = 10'b1010101100;
mem2[9365] = 10'b1010101101;
mem2[9366] = 10'b1010101101;
mem2[9367] = 10'b1010101101;
mem2[9368] = 10'b1010101101;
mem2[9369] = 10'b1010101101;
mem2[9370] = 10'b1010101101;
mem2[9371] = 10'b1010101101;
mem2[9372] = 10'b1010101101;
mem2[9373] = 10'b1010101101;
mem2[9374] = 10'b1010101101;
mem2[9375] = 10'b1010101110;
mem2[9376] = 10'b1010101110;
mem2[9377] = 10'b1010101110;
mem2[9378] = 10'b1010101110;
mem2[9379] = 10'b1010101110;
mem2[9380] = 10'b1010101110;
mem2[9381] = 10'b1010101110;
mem2[9382] = 10'b1010101110;
mem2[9383] = 10'b1010101110;
mem2[9384] = 10'b1010101110;
mem2[9385] = 10'b1010101111;
mem2[9386] = 10'b1010101111;
mem2[9387] = 10'b1010101111;
mem2[9388] = 10'b1010101111;
mem2[9389] = 10'b1010101111;
mem2[9390] = 10'b1010101111;
mem2[9391] = 10'b1010101111;
mem2[9392] = 10'b1010101111;
mem2[9393] = 10'b1010101111;
mem2[9394] = 10'b1010101111;
mem2[9395] = 10'b1010101111;
mem2[9396] = 10'b1010110000;
mem2[9397] = 10'b1010110000;
mem2[9398] = 10'b1010110000;
mem2[9399] = 10'b1010110000;
mem2[9400] = 10'b1010110000;
mem2[9401] = 10'b1010110000;
mem2[9402] = 10'b1010110000;
mem2[9403] = 10'b1010110000;
mem2[9404] = 10'b1010110000;
mem2[9405] = 10'b1010110000;
mem2[9406] = 10'b1010110001;
mem2[9407] = 10'b1010110001;
mem2[9408] = 10'b1010110001;
mem2[9409] = 10'b1010110001;
mem2[9410] = 10'b1010110001;
mem2[9411] = 10'b1010110001;
mem2[9412] = 10'b1010110001;
mem2[9413] = 10'b1010110001;
mem2[9414] = 10'b1010110001;
mem2[9415] = 10'b1010110001;
mem2[9416] = 10'b1010110010;
mem2[9417] = 10'b1010110010;
mem2[9418] = 10'b1010110010;
mem2[9419] = 10'b1010110010;
mem2[9420] = 10'b1010110010;
mem2[9421] = 10'b1010110010;
mem2[9422] = 10'b1010110010;
mem2[9423] = 10'b1010110010;
mem2[9424] = 10'b1010110010;
mem2[9425] = 10'b1010110010;
mem2[9426] = 10'b1010110011;
mem2[9427] = 10'b1010110011;
mem2[9428] = 10'b1010110011;
mem2[9429] = 10'b1010110011;
mem2[9430] = 10'b1010110011;
mem2[9431] = 10'b1010110011;
mem2[9432] = 10'b1010110011;
mem2[9433] = 10'b1010110011;
mem2[9434] = 10'b1010110011;
mem2[9435] = 10'b1010110011;
mem2[9436] = 10'b1010110100;
mem2[9437] = 10'b1010110100;
mem2[9438] = 10'b1010110100;
mem2[9439] = 10'b1010110100;
mem2[9440] = 10'b1010110100;
mem2[9441] = 10'b1010110100;
mem2[9442] = 10'b1010110100;
mem2[9443] = 10'b1010110100;
mem2[9444] = 10'b1010110100;
mem2[9445] = 10'b1010110100;
mem2[9446] = 10'b1010110100;
mem2[9447] = 10'b1010110101;
mem2[9448] = 10'b1010110101;
mem2[9449] = 10'b1010110101;
mem2[9450] = 10'b1010110101;
mem2[9451] = 10'b1010110101;
mem2[9452] = 10'b1010110101;
mem2[9453] = 10'b1010110101;
mem2[9454] = 10'b1010110101;
mem2[9455] = 10'b1010110101;
mem2[9456] = 10'b1010110101;
mem2[9457] = 10'b1010110110;
mem2[9458] = 10'b1010110110;
mem2[9459] = 10'b1010110110;
mem2[9460] = 10'b1010110110;
mem2[9461] = 10'b1010110110;
mem2[9462] = 10'b1010110110;
mem2[9463] = 10'b1010110110;
mem2[9464] = 10'b1010110110;
mem2[9465] = 10'b1010110110;
mem2[9466] = 10'b1010110110;
mem2[9467] = 10'b1010110111;
mem2[9468] = 10'b1010110111;
mem2[9469] = 10'b1010110111;
mem2[9470] = 10'b1010110111;
mem2[9471] = 10'b1010110111;
mem2[9472] = 10'b1010110111;
mem2[9473] = 10'b1010110111;
mem2[9474] = 10'b1010110111;
mem2[9475] = 10'b1010110111;
mem2[9476] = 10'b1010110111;
mem2[9477] = 10'b1010111000;
mem2[9478] = 10'b1010111000;
mem2[9479] = 10'b1010111000;
mem2[9480] = 10'b1010111000;
mem2[9481] = 10'b1010111000;
mem2[9482] = 10'b1010111000;
mem2[9483] = 10'b1010111000;
mem2[9484] = 10'b1010111000;
mem2[9485] = 10'b1010111000;
mem2[9486] = 10'b1010111000;
mem2[9487] = 10'b1010111001;
mem2[9488] = 10'b1010111001;
mem2[9489] = 10'b1010111001;
mem2[9490] = 10'b1010111001;
mem2[9491] = 10'b1010111001;
mem2[9492] = 10'b1010111001;
mem2[9493] = 10'b1010111001;
mem2[9494] = 10'b1010111001;
mem2[9495] = 10'b1010111001;
mem2[9496] = 10'b1010111001;
mem2[9497] = 10'b1010111001;
mem2[9498] = 10'b1010111010;
mem2[9499] = 10'b1010111010;
mem2[9500] = 10'b1010111010;
mem2[9501] = 10'b1010111010;
mem2[9502] = 10'b1010111010;
mem2[9503] = 10'b1010111010;
mem2[9504] = 10'b1010111010;
mem2[9505] = 10'b1010111010;
mem2[9506] = 10'b1010111010;
mem2[9507] = 10'b1010111010;
mem2[9508] = 10'b1010111011;
mem2[9509] = 10'b1010111011;
mem2[9510] = 10'b1010111011;
mem2[9511] = 10'b1010111011;
mem2[9512] = 10'b1010111011;
mem2[9513] = 10'b1010111011;
mem2[9514] = 10'b1010111011;
mem2[9515] = 10'b1010111011;
mem2[9516] = 10'b1010111011;
mem2[9517] = 10'b1010111011;
mem2[9518] = 10'b1010111100;
mem2[9519] = 10'b1010111100;
mem2[9520] = 10'b1010111100;
mem2[9521] = 10'b1010111100;
mem2[9522] = 10'b1010111100;
mem2[9523] = 10'b1010111100;
mem2[9524] = 10'b1010111100;
mem2[9525] = 10'b1010111100;
mem2[9526] = 10'b1010111100;
mem2[9527] = 10'b1010111100;
mem2[9528] = 10'b1010111101;
mem2[9529] = 10'b1010111101;
mem2[9530] = 10'b1010111101;
mem2[9531] = 10'b1010111101;
mem2[9532] = 10'b1010111101;
mem2[9533] = 10'b1010111101;
mem2[9534] = 10'b1010111101;
mem2[9535] = 10'b1010111101;
mem2[9536] = 10'b1010111101;
mem2[9537] = 10'b1010111101;
mem2[9538] = 10'b1010111101;
mem2[9539] = 10'b1010111110;
mem2[9540] = 10'b1010111110;
mem2[9541] = 10'b1010111110;
mem2[9542] = 10'b1010111110;
mem2[9543] = 10'b1010111110;
mem2[9544] = 10'b1010111110;
mem2[9545] = 10'b1010111110;
mem2[9546] = 10'b1010111110;
mem2[9547] = 10'b1010111110;
mem2[9548] = 10'b1010111110;
mem2[9549] = 10'b1010111111;
mem2[9550] = 10'b1010111111;
mem2[9551] = 10'b1010111111;
mem2[9552] = 10'b1010111111;
mem2[9553] = 10'b1010111111;
mem2[9554] = 10'b1010111111;
mem2[9555] = 10'b1010111111;
mem2[9556] = 10'b1010111111;
mem2[9557] = 10'b1010111111;
mem2[9558] = 10'b1010111111;
mem2[9559] = 10'b1011000000;
mem2[9560] = 10'b1011000000;
mem2[9561] = 10'b1011000000;
mem2[9562] = 10'b1011000000;
mem2[9563] = 10'b1011000000;
mem2[9564] = 10'b1011000000;
mem2[9565] = 10'b1011000000;
mem2[9566] = 10'b1011000000;
mem2[9567] = 10'b1011000000;
mem2[9568] = 10'b1011000000;
mem2[9569] = 10'b1011000000;
mem2[9570] = 10'b1011000001;
mem2[9571] = 10'b1011000001;
mem2[9572] = 10'b1011000001;
mem2[9573] = 10'b1011000001;
mem2[9574] = 10'b1011000001;
mem2[9575] = 10'b1011000001;
mem2[9576] = 10'b1011000001;
mem2[9577] = 10'b1011000001;
mem2[9578] = 10'b1011000001;
mem2[9579] = 10'b1011000001;
mem2[9580] = 10'b1011000010;
mem2[9581] = 10'b1011000010;
mem2[9582] = 10'b1011000010;
mem2[9583] = 10'b1011000010;
mem2[9584] = 10'b1011000010;
mem2[9585] = 10'b1011000010;
mem2[9586] = 10'b1011000010;
mem2[9587] = 10'b1011000010;
mem2[9588] = 10'b1011000010;
mem2[9589] = 10'b1011000010;
mem2[9590] = 10'b1011000011;
mem2[9591] = 10'b1011000011;
mem2[9592] = 10'b1011000011;
mem2[9593] = 10'b1011000011;
mem2[9594] = 10'b1011000011;
mem2[9595] = 10'b1011000011;
mem2[9596] = 10'b1011000011;
mem2[9597] = 10'b1011000011;
mem2[9598] = 10'b1011000011;
mem2[9599] = 10'b1011000011;
mem2[9600] = 10'b1011000011;
mem2[9601] = 10'b1011000100;
mem2[9602] = 10'b1011000100;
mem2[9603] = 10'b1011000100;
mem2[9604] = 10'b1011000100;
mem2[9605] = 10'b1011000100;
mem2[9606] = 10'b1011000100;
mem2[9607] = 10'b1011000100;
mem2[9608] = 10'b1011000100;
mem2[9609] = 10'b1011000100;
mem2[9610] = 10'b1011000100;
mem2[9611] = 10'b1011000101;
mem2[9612] = 10'b1011000101;
mem2[9613] = 10'b1011000101;
mem2[9614] = 10'b1011000101;
mem2[9615] = 10'b1011000101;
mem2[9616] = 10'b1011000101;
mem2[9617] = 10'b1011000101;
mem2[9618] = 10'b1011000101;
mem2[9619] = 10'b1011000101;
mem2[9620] = 10'b1011000101;
mem2[9621] = 10'b1011000110;
mem2[9622] = 10'b1011000110;
mem2[9623] = 10'b1011000110;
mem2[9624] = 10'b1011000110;
mem2[9625] = 10'b1011000110;
mem2[9626] = 10'b1011000110;
mem2[9627] = 10'b1011000110;
mem2[9628] = 10'b1011000110;
mem2[9629] = 10'b1011000110;
mem2[9630] = 10'b1011000110;
mem2[9631] = 10'b1011000110;
mem2[9632] = 10'b1011000111;
mem2[9633] = 10'b1011000111;
mem2[9634] = 10'b1011000111;
mem2[9635] = 10'b1011000111;
mem2[9636] = 10'b1011000111;
mem2[9637] = 10'b1011000111;
mem2[9638] = 10'b1011000111;
mem2[9639] = 10'b1011000111;
mem2[9640] = 10'b1011000111;
mem2[9641] = 10'b1011000111;
mem2[9642] = 10'b1011001000;
mem2[9643] = 10'b1011001000;
mem2[9644] = 10'b1011001000;
mem2[9645] = 10'b1011001000;
mem2[9646] = 10'b1011001000;
mem2[9647] = 10'b1011001000;
mem2[9648] = 10'b1011001000;
mem2[9649] = 10'b1011001000;
mem2[9650] = 10'b1011001000;
mem2[9651] = 10'b1011001000;
mem2[9652] = 10'b1011001001;
mem2[9653] = 10'b1011001001;
mem2[9654] = 10'b1011001001;
mem2[9655] = 10'b1011001001;
mem2[9656] = 10'b1011001001;
mem2[9657] = 10'b1011001001;
mem2[9658] = 10'b1011001001;
mem2[9659] = 10'b1011001001;
mem2[9660] = 10'b1011001001;
mem2[9661] = 10'b1011001001;
mem2[9662] = 10'b1011001001;
mem2[9663] = 10'b1011001010;
mem2[9664] = 10'b1011001010;
mem2[9665] = 10'b1011001010;
mem2[9666] = 10'b1011001010;
mem2[9667] = 10'b1011001010;
mem2[9668] = 10'b1011001010;
mem2[9669] = 10'b1011001010;
mem2[9670] = 10'b1011001010;
mem2[9671] = 10'b1011001010;
mem2[9672] = 10'b1011001010;
mem2[9673] = 10'b1011001011;
mem2[9674] = 10'b1011001011;
mem2[9675] = 10'b1011001011;
mem2[9676] = 10'b1011001011;
mem2[9677] = 10'b1011001011;
mem2[9678] = 10'b1011001011;
mem2[9679] = 10'b1011001011;
mem2[9680] = 10'b1011001011;
mem2[9681] = 10'b1011001011;
mem2[9682] = 10'b1011001011;
mem2[9683] = 10'b1011001011;
mem2[9684] = 10'b1011001100;
mem2[9685] = 10'b1011001100;
mem2[9686] = 10'b1011001100;
mem2[9687] = 10'b1011001100;
mem2[9688] = 10'b1011001100;
mem2[9689] = 10'b1011001100;
mem2[9690] = 10'b1011001100;
mem2[9691] = 10'b1011001100;
mem2[9692] = 10'b1011001100;
mem2[9693] = 10'b1011001100;
mem2[9694] = 10'b1011001101;
mem2[9695] = 10'b1011001101;
mem2[9696] = 10'b1011001101;
mem2[9697] = 10'b1011001101;
mem2[9698] = 10'b1011001101;
mem2[9699] = 10'b1011001101;
mem2[9700] = 10'b1011001101;
mem2[9701] = 10'b1011001101;
mem2[9702] = 10'b1011001101;
mem2[9703] = 10'b1011001101;
mem2[9704] = 10'b1011001110;
mem2[9705] = 10'b1011001110;
mem2[9706] = 10'b1011001110;
mem2[9707] = 10'b1011001110;
mem2[9708] = 10'b1011001110;
mem2[9709] = 10'b1011001110;
mem2[9710] = 10'b1011001110;
mem2[9711] = 10'b1011001110;
mem2[9712] = 10'b1011001110;
mem2[9713] = 10'b1011001110;
mem2[9714] = 10'b1011001110;
mem2[9715] = 10'b1011001111;
mem2[9716] = 10'b1011001111;
mem2[9717] = 10'b1011001111;
mem2[9718] = 10'b1011001111;
mem2[9719] = 10'b1011001111;
mem2[9720] = 10'b1011001111;
mem2[9721] = 10'b1011001111;
mem2[9722] = 10'b1011001111;
mem2[9723] = 10'b1011001111;
mem2[9724] = 10'b1011001111;
mem2[9725] = 10'b1011010000;
mem2[9726] = 10'b1011010000;
mem2[9727] = 10'b1011010000;
mem2[9728] = 10'b1011010000;
mem2[9729] = 10'b1011010000;
mem2[9730] = 10'b1011010000;
mem2[9731] = 10'b1011010000;
mem2[9732] = 10'b1011010000;
mem2[9733] = 10'b1011010000;
mem2[9734] = 10'b1011010000;
mem2[9735] = 10'b1011010000;
mem2[9736] = 10'b1011010001;
mem2[9737] = 10'b1011010001;
mem2[9738] = 10'b1011010001;
mem2[9739] = 10'b1011010001;
mem2[9740] = 10'b1011010001;
mem2[9741] = 10'b1011010001;
mem2[9742] = 10'b1011010001;
mem2[9743] = 10'b1011010001;
mem2[9744] = 10'b1011010001;
mem2[9745] = 10'b1011010001;
mem2[9746] = 10'b1011010010;
mem2[9747] = 10'b1011010010;
mem2[9748] = 10'b1011010010;
mem2[9749] = 10'b1011010010;
mem2[9750] = 10'b1011010010;
mem2[9751] = 10'b1011010010;
mem2[9752] = 10'b1011010010;
mem2[9753] = 10'b1011010010;
mem2[9754] = 10'b1011010010;
mem2[9755] = 10'b1011010010;
mem2[9756] = 10'b1011010010;
mem2[9757] = 10'b1011010011;
mem2[9758] = 10'b1011010011;
mem2[9759] = 10'b1011010011;
mem2[9760] = 10'b1011010011;
mem2[9761] = 10'b1011010011;
mem2[9762] = 10'b1011010011;
mem2[9763] = 10'b1011010011;
mem2[9764] = 10'b1011010011;
mem2[9765] = 10'b1011010011;
mem2[9766] = 10'b1011010011;
mem2[9767] = 10'b1011010100;
mem2[9768] = 10'b1011010100;
mem2[9769] = 10'b1011010100;
mem2[9770] = 10'b1011010100;
mem2[9771] = 10'b1011010100;
mem2[9772] = 10'b1011010100;
mem2[9773] = 10'b1011010100;
mem2[9774] = 10'b1011010100;
mem2[9775] = 10'b1011010100;
mem2[9776] = 10'b1011010100;
mem2[9777] = 10'b1011010100;
mem2[9778] = 10'b1011010101;
mem2[9779] = 10'b1011010101;
mem2[9780] = 10'b1011010101;
mem2[9781] = 10'b1011010101;
mem2[9782] = 10'b1011010101;
mem2[9783] = 10'b1011010101;
mem2[9784] = 10'b1011010101;
mem2[9785] = 10'b1011010101;
mem2[9786] = 10'b1011010101;
mem2[9787] = 10'b1011010101;
mem2[9788] = 10'b1011010110;
mem2[9789] = 10'b1011010110;
mem2[9790] = 10'b1011010110;
mem2[9791] = 10'b1011010110;
mem2[9792] = 10'b1011010110;
mem2[9793] = 10'b1011010110;
mem2[9794] = 10'b1011010110;
mem2[9795] = 10'b1011010110;
mem2[9796] = 10'b1011010110;
mem2[9797] = 10'b1011010110;
mem2[9798] = 10'b1011010110;
mem2[9799] = 10'b1011010111;
mem2[9800] = 10'b1011010111;
mem2[9801] = 10'b1011010111;
mem2[9802] = 10'b1011010111;
mem2[9803] = 10'b1011010111;
mem2[9804] = 10'b1011010111;
mem2[9805] = 10'b1011010111;
mem2[9806] = 10'b1011010111;
mem2[9807] = 10'b1011010111;
mem2[9808] = 10'b1011010111;
mem2[9809] = 10'b1011011000;
mem2[9810] = 10'b1011011000;
mem2[9811] = 10'b1011011000;
mem2[9812] = 10'b1011011000;
mem2[9813] = 10'b1011011000;
mem2[9814] = 10'b1011011000;
mem2[9815] = 10'b1011011000;
mem2[9816] = 10'b1011011000;
mem2[9817] = 10'b1011011000;
mem2[9818] = 10'b1011011000;
mem2[9819] = 10'b1011011000;
mem2[9820] = 10'b1011011001;
mem2[9821] = 10'b1011011001;
mem2[9822] = 10'b1011011001;
mem2[9823] = 10'b1011011001;
mem2[9824] = 10'b1011011001;
mem2[9825] = 10'b1011011001;
mem2[9826] = 10'b1011011001;
mem2[9827] = 10'b1011011001;
mem2[9828] = 10'b1011011001;
mem2[9829] = 10'b1011011001;
mem2[9830] = 10'b1011011010;
mem2[9831] = 10'b1011011010;
mem2[9832] = 10'b1011011010;
mem2[9833] = 10'b1011011010;
mem2[9834] = 10'b1011011010;
mem2[9835] = 10'b1011011010;
mem2[9836] = 10'b1011011010;
mem2[9837] = 10'b1011011010;
mem2[9838] = 10'b1011011010;
mem2[9839] = 10'b1011011010;
mem2[9840] = 10'b1011011010;
mem2[9841] = 10'b1011011011;
mem2[9842] = 10'b1011011011;
mem2[9843] = 10'b1011011011;
mem2[9844] = 10'b1011011011;
mem2[9845] = 10'b1011011011;
mem2[9846] = 10'b1011011011;
mem2[9847] = 10'b1011011011;
mem2[9848] = 10'b1011011011;
mem2[9849] = 10'b1011011011;
mem2[9850] = 10'b1011011011;
mem2[9851] = 10'b1011011100;
mem2[9852] = 10'b1011011100;
mem2[9853] = 10'b1011011100;
mem2[9854] = 10'b1011011100;
mem2[9855] = 10'b1011011100;
mem2[9856] = 10'b1011011100;
mem2[9857] = 10'b1011011100;
mem2[9858] = 10'b1011011100;
mem2[9859] = 10'b1011011100;
mem2[9860] = 10'b1011011100;
mem2[9861] = 10'b1011011100;
mem2[9862] = 10'b1011011101;
mem2[9863] = 10'b1011011101;
mem2[9864] = 10'b1011011101;
mem2[9865] = 10'b1011011101;
mem2[9866] = 10'b1011011101;
mem2[9867] = 10'b1011011101;
mem2[9868] = 10'b1011011101;
mem2[9869] = 10'b1011011101;
mem2[9870] = 10'b1011011101;
mem2[9871] = 10'b1011011101;
mem2[9872] = 10'b1011011101;
mem2[9873] = 10'b1011011110;
mem2[9874] = 10'b1011011110;
mem2[9875] = 10'b1011011110;
mem2[9876] = 10'b1011011110;
mem2[9877] = 10'b1011011110;
mem2[9878] = 10'b1011011110;
mem2[9879] = 10'b1011011110;
mem2[9880] = 10'b1011011110;
mem2[9881] = 10'b1011011110;
mem2[9882] = 10'b1011011110;
mem2[9883] = 10'b1011011111;
mem2[9884] = 10'b1011011111;
mem2[9885] = 10'b1011011111;
mem2[9886] = 10'b1011011111;
mem2[9887] = 10'b1011011111;
mem2[9888] = 10'b1011011111;
mem2[9889] = 10'b1011011111;
mem2[9890] = 10'b1011011111;
mem2[9891] = 10'b1011011111;
mem2[9892] = 10'b1011011111;
mem2[9893] = 10'b1011011111;
mem2[9894] = 10'b1011100000;
mem2[9895] = 10'b1011100000;
mem2[9896] = 10'b1011100000;
mem2[9897] = 10'b1011100000;
mem2[9898] = 10'b1011100000;
mem2[9899] = 10'b1011100000;
mem2[9900] = 10'b1011100000;
mem2[9901] = 10'b1011100000;
mem2[9902] = 10'b1011100000;
mem2[9903] = 10'b1011100000;
mem2[9904] = 10'b1011100001;
mem2[9905] = 10'b1011100001;
mem2[9906] = 10'b1011100001;
mem2[9907] = 10'b1011100001;
mem2[9908] = 10'b1011100001;
mem2[9909] = 10'b1011100001;
mem2[9910] = 10'b1011100001;
mem2[9911] = 10'b1011100001;
mem2[9912] = 10'b1011100001;
mem2[9913] = 10'b1011100001;
mem2[9914] = 10'b1011100001;
mem2[9915] = 10'b1011100010;
mem2[9916] = 10'b1011100010;
mem2[9917] = 10'b1011100010;
mem2[9918] = 10'b1011100010;
mem2[9919] = 10'b1011100010;
mem2[9920] = 10'b1011100010;
mem2[9921] = 10'b1011100010;
mem2[9922] = 10'b1011100010;
mem2[9923] = 10'b1011100010;
mem2[9924] = 10'b1011100010;
mem2[9925] = 10'b1011100010;
mem2[9926] = 10'b1011100011;
mem2[9927] = 10'b1011100011;
mem2[9928] = 10'b1011100011;
mem2[9929] = 10'b1011100011;
mem2[9930] = 10'b1011100011;
mem2[9931] = 10'b1011100011;
mem2[9932] = 10'b1011100011;
mem2[9933] = 10'b1011100011;
mem2[9934] = 10'b1011100011;
mem2[9935] = 10'b1011100011;
mem2[9936] = 10'b1011100100;
mem2[9937] = 10'b1011100100;
mem2[9938] = 10'b1011100100;
mem2[9939] = 10'b1011100100;
mem2[9940] = 10'b1011100100;
mem2[9941] = 10'b1011100100;
mem2[9942] = 10'b1011100100;
mem2[9943] = 10'b1011100100;
mem2[9944] = 10'b1011100100;
mem2[9945] = 10'b1011100100;
mem2[9946] = 10'b1011100100;
mem2[9947] = 10'b1011100101;
mem2[9948] = 10'b1011100101;
mem2[9949] = 10'b1011100101;
mem2[9950] = 10'b1011100101;
mem2[9951] = 10'b1011100101;
mem2[9952] = 10'b1011100101;
mem2[9953] = 10'b1011100101;
mem2[9954] = 10'b1011100101;
mem2[9955] = 10'b1011100101;
mem2[9956] = 10'b1011100101;
mem2[9957] = 10'b1011100101;
mem2[9958] = 10'b1011100110;
mem2[9959] = 10'b1011100110;
mem2[9960] = 10'b1011100110;
mem2[9961] = 10'b1011100110;
mem2[9962] = 10'b1011100110;
mem2[9963] = 10'b1011100110;
mem2[9964] = 10'b1011100110;
mem2[9965] = 10'b1011100110;
mem2[9966] = 10'b1011100110;
mem2[9967] = 10'b1011100110;
mem2[9968] = 10'b1011100111;
mem2[9969] = 10'b1011100111;
mem2[9970] = 10'b1011100111;
mem2[9971] = 10'b1011100111;
mem2[9972] = 10'b1011100111;
mem2[9973] = 10'b1011100111;
mem2[9974] = 10'b1011100111;
mem2[9975] = 10'b1011100111;
mem2[9976] = 10'b1011100111;
mem2[9977] = 10'b1011100111;
mem2[9978] = 10'b1011100111;
mem2[9979] = 10'b1011101000;
mem2[9980] = 10'b1011101000;
mem2[9981] = 10'b1011101000;
mem2[9982] = 10'b1011101000;
mem2[9983] = 10'b1011101000;
mem2[9984] = 10'b1011101000;
mem2[9985] = 10'b1011101000;
mem2[9986] = 10'b1011101000;
mem2[9987] = 10'b1011101000;
mem2[9988] = 10'b1011101000;
mem2[9989] = 10'b1011101000;
mem2[9990] = 10'b1011101001;
mem2[9991] = 10'b1011101001;
mem2[9992] = 10'b1011101001;
mem2[9993] = 10'b1011101001;
mem2[9994] = 10'b1011101001;
mem2[9995] = 10'b1011101001;
mem2[9996] = 10'b1011101001;
mem2[9997] = 10'b1011101001;
mem2[9998] = 10'b1011101001;
mem2[9999] = 10'b1011101001;
mem2[10000] = 10'b1011101001;
mem2[10001] = 10'b1011101010;
mem2[10002] = 10'b1011101010;
mem2[10003] = 10'b1011101010;
mem2[10004] = 10'b1011101010;
mem2[10005] = 10'b1011101010;
mem2[10006] = 10'b1011101010;
mem2[10007] = 10'b1011101010;
mem2[10008] = 10'b1011101010;
mem2[10009] = 10'b1011101010;
mem2[10010] = 10'b1011101010;
mem2[10011] = 10'b1011101011;
mem2[10012] = 10'b1011101011;
mem2[10013] = 10'b1011101011;
mem2[10014] = 10'b1011101011;
mem2[10015] = 10'b1011101011;
mem2[10016] = 10'b1011101011;
mem2[10017] = 10'b1011101011;
mem2[10018] = 10'b1011101011;
mem2[10019] = 10'b1011101011;
mem2[10020] = 10'b1011101011;
mem2[10021] = 10'b1011101011;
mem2[10022] = 10'b1011101100;
mem2[10023] = 10'b1011101100;
mem2[10024] = 10'b1011101100;
mem2[10025] = 10'b1011101100;
mem2[10026] = 10'b1011101100;
mem2[10027] = 10'b1011101100;
mem2[10028] = 10'b1011101100;
mem2[10029] = 10'b1011101100;
mem2[10030] = 10'b1011101100;
mem2[10031] = 10'b1011101100;
mem2[10032] = 10'b1011101100;
mem2[10033] = 10'b1011101101;
mem2[10034] = 10'b1011101101;
mem2[10035] = 10'b1011101101;
mem2[10036] = 10'b1011101101;
mem2[10037] = 10'b1011101101;
mem2[10038] = 10'b1011101101;
mem2[10039] = 10'b1011101101;
mem2[10040] = 10'b1011101101;
mem2[10041] = 10'b1011101101;
mem2[10042] = 10'b1011101101;
mem2[10043] = 10'b1011101101;
mem2[10044] = 10'b1011101110;
mem2[10045] = 10'b1011101110;
mem2[10046] = 10'b1011101110;
mem2[10047] = 10'b1011101110;
mem2[10048] = 10'b1011101110;
mem2[10049] = 10'b1011101110;
mem2[10050] = 10'b1011101110;
mem2[10051] = 10'b1011101110;
mem2[10052] = 10'b1011101110;
mem2[10053] = 10'b1011101110;
mem2[10054] = 10'b1011101111;
mem2[10055] = 10'b1011101111;
mem2[10056] = 10'b1011101111;
mem2[10057] = 10'b1011101111;
mem2[10058] = 10'b1011101111;
mem2[10059] = 10'b1011101111;
mem2[10060] = 10'b1011101111;
mem2[10061] = 10'b1011101111;
mem2[10062] = 10'b1011101111;
mem2[10063] = 10'b1011101111;
mem2[10064] = 10'b1011101111;
mem2[10065] = 10'b1011110000;
mem2[10066] = 10'b1011110000;
mem2[10067] = 10'b1011110000;
mem2[10068] = 10'b1011110000;
mem2[10069] = 10'b1011110000;
mem2[10070] = 10'b1011110000;
mem2[10071] = 10'b1011110000;
mem2[10072] = 10'b1011110000;
mem2[10073] = 10'b1011110000;
mem2[10074] = 10'b1011110000;
mem2[10075] = 10'b1011110000;
mem2[10076] = 10'b1011110001;
mem2[10077] = 10'b1011110001;
mem2[10078] = 10'b1011110001;
mem2[10079] = 10'b1011110001;
mem2[10080] = 10'b1011110001;
mem2[10081] = 10'b1011110001;
mem2[10082] = 10'b1011110001;
mem2[10083] = 10'b1011110001;
mem2[10084] = 10'b1011110001;
mem2[10085] = 10'b1011110001;
mem2[10086] = 10'b1011110001;
mem2[10087] = 10'b1011110010;
mem2[10088] = 10'b1011110010;
mem2[10089] = 10'b1011110010;
mem2[10090] = 10'b1011110010;
mem2[10091] = 10'b1011110010;
mem2[10092] = 10'b1011110010;
mem2[10093] = 10'b1011110010;
mem2[10094] = 10'b1011110010;
mem2[10095] = 10'b1011110010;
mem2[10096] = 10'b1011110010;
mem2[10097] = 10'b1011110010;
mem2[10098] = 10'b1011110011;
mem2[10099] = 10'b1011110011;
mem2[10100] = 10'b1011110011;
mem2[10101] = 10'b1011110011;
mem2[10102] = 10'b1011110011;
mem2[10103] = 10'b1011110011;
mem2[10104] = 10'b1011110011;
mem2[10105] = 10'b1011110011;
mem2[10106] = 10'b1011110011;
mem2[10107] = 10'b1011110011;
mem2[10108] = 10'b1011110011;
mem2[10109] = 10'b1011110100;
mem2[10110] = 10'b1011110100;
mem2[10111] = 10'b1011110100;
mem2[10112] = 10'b1011110100;
mem2[10113] = 10'b1011110100;
mem2[10114] = 10'b1011110100;
mem2[10115] = 10'b1011110100;
mem2[10116] = 10'b1011110100;
mem2[10117] = 10'b1011110100;
mem2[10118] = 10'b1011110100;
mem2[10119] = 10'b1011110101;
mem2[10120] = 10'b1011110101;
mem2[10121] = 10'b1011110101;
mem2[10122] = 10'b1011110101;
mem2[10123] = 10'b1011110101;
mem2[10124] = 10'b1011110101;
mem2[10125] = 10'b1011110101;
mem2[10126] = 10'b1011110101;
mem2[10127] = 10'b1011110101;
mem2[10128] = 10'b1011110101;
mem2[10129] = 10'b1011110101;
mem2[10130] = 10'b1011110110;
mem2[10131] = 10'b1011110110;
mem2[10132] = 10'b1011110110;
mem2[10133] = 10'b1011110110;
mem2[10134] = 10'b1011110110;
mem2[10135] = 10'b1011110110;
mem2[10136] = 10'b1011110110;
mem2[10137] = 10'b1011110110;
mem2[10138] = 10'b1011110110;
mem2[10139] = 10'b1011110110;
mem2[10140] = 10'b1011110110;
mem2[10141] = 10'b1011110111;
mem2[10142] = 10'b1011110111;
mem2[10143] = 10'b1011110111;
mem2[10144] = 10'b1011110111;
mem2[10145] = 10'b1011110111;
mem2[10146] = 10'b1011110111;
mem2[10147] = 10'b1011110111;
mem2[10148] = 10'b1011110111;
mem2[10149] = 10'b1011110111;
mem2[10150] = 10'b1011110111;
mem2[10151] = 10'b1011110111;
mem2[10152] = 10'b1011111000;
mem2[10153] = 10'b1011111000;
mem2[10154] = 10'b1011111000;
mem2[10155] = 10'b1011111000;
mem2[10156] = 10'b1011111000;
mem2[10157] = 10'b1011111000;
mem2[10158] = 10'b1011111000;
mem2[10159] = 10'b1011111000;
mem2[10160] = 10'b1011111000;
mem2[10161] = 10'b1011111000;
mem2[10162] = 10'b1011111000;
mem2[10163] = 10'b1011111001;
mem2[10164] = 10'b1011111001;
mem2[10165] = 10'b1011111001;
mem2[10166] = 10'b1011111001;
mem2[10167] = 10'b1011111001;
mem2[10168] = 10'b1011111001;
mem2[10169] = 10'b1011111001;
mem2[10170] = 10'b1011111001;
mem2[10171] = 10'b1011111001;
mem2[10172] = 10'b1011111001;
mem2[10173] = 10'b1011111001;
mem2[10174] = 10'b1011111010;
mem2[10175] = 10'b1011111010;
mem2[10176] = 10'b1011111010;
mem2[10177] = 10'b1011111010;
mem2[10178] = 10'b1011111010;
mem2[10179] = 10'b1011111010;
mem2[10180] = 10'b1011111010;
mem2[10181] = 10'b1011111010;
mem2[10182] = 10'b1011111010;
mem2[10183] = 10'b1011111010;
mem2[10184] = 10'b1011111010;
mem2[10185] = 10'b1011111011;
mem2[10186] = 10'b1011111011;
mem2[10187] = 10'b1011111011;
mem2[10188] = 10'b1011111011;
mem2[10189] = 10'b1011111011;
mem2[10190] = 10'b1011111011;
mem2[10191] = 10'b1011111011;
mem2[10192] = 10'b1011111011;
mem2[10193] = 10'b1011111011;
mem2[10194] = 10'b1011111011;
mem2[10195] = 10'b1011111011;
mem2[10196] = 10'b1011111100;
mem2[10197] = 10'b1011111100;
mem2[10198] = 10'b1011111100;
mem2[10199] = 10'b1011111100;
mem2[10200] = 10'b1011111100;
mem2[10201] = 10'b1011111100;
mem2[10202] = 10'b1011111100;
mem2[10203] = 10'b1011111100;
mem2[10204] = 10'b1011111100;
mem2[10205] = 10'b1011111100;
mem2[10206] = 10'b1011111100;
mem2[10207] = 10'b1011111101;
mem2[10208] = 10'b1011111101;
mem2[10209] = 10'b1011111101;
mem2[10210] = 10'b1011111101;
mem2[10211] = 10'b1011111101;
mem2[10212] = 10'b1011111101;
mem2[10213] = 10'b1011111101;
mem2[10214] = 10'b1011111101;
mem2[10215] = 10'b1011111101;
mem2[10216] = 10'b1011111101;
mem2[10217] = 10'b1011111101;
mem2[10218] = 10'b1011111110;
mem2[10219] = 10'b1011111110;
mem2[10220] = 10'b1011111110;
mem2[10221] = 10'b1011111110;
mem2[10222] = 10'b1011111110;
mem2[10223] = 10'b1011111110;
mem2[10224] = 10'b1011111110;
mem2[10225] = 10'b1011111110;
mem2[10226] = 10'b1011111110;
mem2[10227] = 10'b1011111110;
mem2[10228] = 10'b1011111110;
mem2[10229] = 10'b1011111111;
mem2[10230] = 10'b1011111111;
mem2[10231] = 10'b1011111111;
mem2[10232] = 10'b1011111111;
mem2[10233] = 10'b1011111111;
mem2[10234] = 10'b1011111111;
mem2[10235] = 10'b1011111111;
mem2[10236] = 10'b1011111111;
mem2[10237] = 10'b1011111111;
mem2[10238] = 10'b1011111111;
mem2[10239] = 10'b1011111111;
mem2[10240] = 10'b1100000000;
mem2[10241] = 10'b1100000000;
mem2[10242] = 10'b1100000000;
mem2[10243] = 10'b1100000000;
mem2[10244] = 10'b1100000000;
mem2[10245] = 10'b1100000000;
mem2[10246] = 10'b1100000000;
mem2[10247] = 10'b1100000000;
mem2[10248] = 10'b1100000000;
mem2[10249] = 10'b1100000000;
mem2[10250] = 10'b1100000000;
mem2[10251] = 10'b1100000001;
mem2[10252] = 10'b1100000001;
mem2[10253] = 10'b1100000001;
mem2[10254] = 10'b1100000001;
mem2[10255] = 10'b1100000001;
mem2[10256] = 10'b1100000001;
mem2[10257] = 10'b1100000001;
mem2[10258] = 10'b1100000001;
mem2[10259] = 10'b1100000001;
mem2[10260] = 10'b1100000001;
mem2[10261] = 10'b1100000001;
mem2[10262] = 10'b1100000010;
mem2[10263] = 10'b1100000010;
mem2[10264] = 10'b1100000010;
mem2[10265] = 10'b1100000010;
mem2[10266] = 10'b1100000010;
mem2[10267] = 10'b1100000010;
mem2[10268] = 10'b1100000010;
mem2[10269] = 10'b1100000010;
mem2[10270] = 10'b1100000010;
mem2[10271] = 10'b1100000010;
mem2[10272] = 10'b1100000010;
mem2[10273] = 10'b1100000011;
mem2[10274] = 10'b1100000011;
mem2[10275] = 10'b1100000011;
mem2[10276] = 10'b1100000011;
mem2[10277] = 10'b1100000011;
mem2[10278] = 10'b1100000011;
mem2[10279] = 10'b1100000011;
mem2[10280] = 10'b1100000011;
mem2[10281] = 10'b1100000011;
mem2[10282] = 10'b1100000011;
mem2[10283] = 10'b1100000011;
mem2[10284] = 10'b1100000100;
mem2[10285] = 10'b1100000100;
mem2[10286] = 10'b1100000100;
mem2[10287] = 10'b1100000100;
mem2[10288] = 10'b1100000100;
mem2[10289] = 10'b1100000100;
mem2[10290] = 10'b1100000100;
mem2[10291] = 10'b1100000100;
mem2[10292] = 10'b1100000100;
mem2[10293] = 10'b1100000100;
mem2[10294] = 10'b1100000100;
mem2[10295] = 10'b1100000101;
mem2[10296] = 10'b1100000101;
mem2[10297] = 10'b1100000101;
mem2[10298] = 10'b1100000101;
mem2[10299] = 10'b1100000101;
mem2[10300] = 10'b1100000101;
mem2[10301] = 10'b1100000101;
mem2[10302] = 10'b1100000101;
mem2[10303] = 10'b1100000101;
mem2[10304] = 10'b1100000101;
mem2[10305] = 10'b1100000101;
mem2[10306] = 10'b1100000110;
mem2[10307] = 10'b1100000110;
mem2[10308] = 10'b1100000110;
mem2[10309] = 10'b1100000110;
mem2[10310] = 10'b1100000110;
mem2[10311] = 10'b1100000110;
mem2[10312] = 10'b1100000110;
mem2[10313] = 10'b1100000110;
mem2[10314] = 10'b1100000110;
mem2[10315] = 10'b1100000110;
mem2[10316] = 10'b1100000110;
mem2[10317] = 10'b1100000111;
mem2[10318] = 10'b1100000111;
mem2[10319] = 10'b1100000111;
mem2[10320] = 10'b1100000111;
mem2[10321] = 10'b1100000111;
mem2[10322] = 10'b1100000111;
mem2[10323] = 10'b1100000111;
mem2[10324] = 10'b1100000111;
mem2[10325] = 10'b1100000111;
mem2[10326] = 10'b1100000111;
mem2[10327] = 10'b1100000111;
mem2[10328] = 10'b1100000111;
mem2[10329] = 10'b1100001000;
mem2[10330] = 10'b1100001000;
mem2[10331] = 10'b1100001000;
mem2[10332] = 10'b1100001000;
mem2[10333] = 10'b1100001000;
mem2[10334] = 10'b1100001000;
mem2[10335] = 10'b1100001000;
mem2[10336] = 10'b1100001000;
mem2[10337] = 10'b1100001000;
mem2[10338] = 10'b1100001000;
mem2[10339] = 10'b1100001000;
mem2[10340] = 10'b1100001001;
mem2[10341] = 10'b1100001001;
mem2[10342] = 10'b1100001001;
mem2[10343] = 10'b1100001001;
mem2[10344] = 10'b1100001001;
mem2[10345] = 10'b1100001001;
mem2[10346] = 10'b1100001001;
mem2[10347] = 10'b1100001001;
mem2[10348] = 10'b1100001001;
mem2[10349] = 10'b1100001001;
mem2[10350] = 10'b1100001001;
mem2[10351] = 10'b1100001010;
mem2[10352] = 10'b1100001010;
mem2[10353] = 10'b1100001010;
mem2[10354] = 10'b1100001010;
mem2[10355] = 10'b1100001010;
mem2[10356] = 10'b1100001010;
mem2[10357] = 10'b1100001010;
mem2[10358] = 10'b1100001010;
mem2[10359] = 10'b1100001010;
mem2[10360] = 10'b1100001010;
mem2[10361] = 10'b1100001010;
mem2[10362] = 10'b1100001011;
mem2[10363] = 10'b1100001011;
mem2[10364] = 10'b1100001011;
mem2[10365] = 10'b1100001011;
mem2[10366] = 10'b1100001011;
mem2[10367] = 10'b1100001011;
mem2[10368] = 10'b1100001011;
mem2[10369] = 10'b1100001011;
mem2[10370] = 10'b1100001011;
mem2[10371] = 10'b1100001011;
mem2[10372] = 10'b1100001011;
mem2[10373] = 10'b1100001100;
mem2[10374] = 10'b1100001100;
mem2[10375] = 10'b1100001100;
mem2[10376] = 10'b1100001100;
mem2[10377] = 10'b1100001100;
mem2[10378] = 10'b1100001100;
mem2[10379] = 10'b1100001100;
mem2[10380] = 10'b1100001100;
mem2[10381] = 10'b1100001100;
mem2[10382] = 10'b1100001100;
mem2[10383] = 10'b1100001100;
mem2[10384] = 10'b1100001100;
mem2[10385] = 10'b1100001101;
mem2[10386] = 10'b1100001101;
mem2[10387] = 10'b1100001101;
mem2[10388] = 10'b1100001101;
mem2[10389] = 10'b1100001101;
mem2[10390] = 10'b1100001101;
mem2[10391] = 10'b1100001101;
mem2[10392] = 10'b1100001101;
mem2[10393] = 10'b1100001101;
mem2[10394] = 10'b1100001101;
mem2[10395] = 10'b1100001101;
mem2[10396] = 10'b1100001110;
mem2[10397] = 10'b1100001110;
mem2[10398] = 10'b1100001110;
mem2[10399] = 10'b1100001110;
mem2[10400] = 10'b1100001110;
mem2[10401] = 10'b1100001110;
mem2[10402] = 10'b1100001110;
mem2[10403] = 10'b1100001110;
mem2[10404] = 10'b1100001110;
mem2[10405] = 10'b1100001110;
mem2[10406] = 10'b1100001110;
mem2[10407] = 10'b1100001111;
mem2[10408] = 10'b1100001111;
mem2[10409] = 10'b1100001111;
mem2[10410] = 10'b1100001111;
mem2[10411] = 10'b1100001111;
mem2[10412] = 10'b1100001111;
mem2[10413] = 10'b1100001111;
mem2[10414] = 10'b1100001111;
mem2[10415] = 10'b1100001111;
mem2[10416] = 10'b1100001111;
mem2[10417] = 10'b1100001111;
mem2[10418] = 10'b1100010000;
mem2[10419] = 10'b1100010000;
mem2[10420] = 10'b1100010000;
mem2[10421] = 10'b1100010000;
mem2[10422] = 10'b1100010000;
mem2[10423] = 10'b1100010000;
mem2[10424] = 10'b1100010000;
mem2[10425] = 10'b1100010000;
mem2[10426] = 10'b1100010000;
mem2[10427] = 10'b1100010000;
mem2[10428] = 10'b1100010000;
mem2[10429] = 10'b1100010000;
mem2[10430] = 10'b1100010001;
mem2[10431] = 10'b1100010001;
mem2[10432] = 10'b1100010001;
mem2[10433] = 10'b1100010001;
mem2[10434] = 10'b1100010001;
mem2[10435] = 10'b1100010001;
mem2[10436] = 10'b1100010001;
mem2[10437] = 10'b1100010001;
mem2[10438] = 10'b1100010001;
mem2[10439] = 10'b1100010001;
mem2[10440] = 10'b1100010001;
mem2[10441] = 10'b1100010010;
mem2[10442] = 10'b1100010010;
mem2[10443] = 10'b1100010010;
mem2[10444] = 10'b1100010010;
mem2[10445] = 10'b1100010010;
mem2[10446] = 10'b1100010010;
mem2[10447] = 10'b1100010010;
mem2[10448] = 10'b1100010010;
mem2[10449] = 10'b1100010010;
mem2[10450] = 10'b1100010010;
mem2[10451] = 10'b1100010010;
mem2[10452] = 10'b1100010011;
mem2[10453] = 10'b1100010011;
mem2[10454] = 10'b1100010011;
mem2[10455] = 10'b1100010011;
mem2[10456] = 10'b1100010011;
mem2[10457] = 10'b1100010011;
mem2[10458] = 10'b1100010011;
mem2[10459] = 10'b1100010011;
mem2[10460] = 10'b1100010011;
mem2[10461] = 10'b1100010011;
mem2[10462] = 10'b1100010011;
mem2[10463] = 10'b1100010100;
mem2[10464] = 10'b1100010100;
mem2[10465] = 10'b1100010100;
mem2[10466] = 10'b1100010100;
mem2[10467] = 10'b1100010100;
mem2[10468] = 10'b1100010100;
mem2[10469] = 10'b1100010100;
mem2[10470] = 10'b1100010100;
mem2[10471] = 10'b1100010100;
mem2[10472] = 10'b1100010100;
mem2[10473] = 10'b1100010100;
mem2[10474] = 10'b1100010100;
mem2[10475] = 10'b1100010101;
mem2[10476] = 10'b1100010101;
mem2[10477] = 10'b1100010101;
mem2[10478] = 10'b1100010101;
mem2[10479] = 10'b1100010101;
mem2[10480] = 10'b1100010101;
mem2[10481] = 10'b1100010101;
mem2[10482] = 10'b1100010101;
mem2[10483] = 10'b1100010101;
mem2[10484] = 10'b1100010101;
mem2[10485] = 10'b1100010101;
mem2[10486] = 10'b1100010110;
mem2[10487] = 10'b1100010110;
mem2[10488] = 10'b1100010110;
mem2[10489] = 10'b1100010110;
mem2[10490] = 10'b1100010110;
mem2[10491] = 10'b1100010110;
mem2[10492] = 10'b1100010110;
mem2[10493] = 10'b1100010110;
mem2[10494] = 10'b1100010110;
mem2[10495] = 10'b1100010110;
mem2[10496] = 10'b1100010110;
mem2[10497] = 10'b1100010110;
mem2[10498] = 10'b1100010111;
mem2[10499] = 10'b1100010111;
mem2[10500] = 10'b1100010111;
mem2[10501] = 10'b1100010111;
mem2[10502] = 10'b1100010111;
mem2[10503] = 10'b1100010111;
mem2[10504] = 10'b1100010111;
mem2[10505] = 10'b1100010111;
mem2[10506] = 10'b1100010111;
mem2[10507] = 10'b1100010111;
mem2[10508] = 10'b1100010111;
mem2[10509] = 10'b1100011000;
mem2[10510] = 10'b1100011000;
mem2[10511] = 10'b1100011000;
mem2[10512] = 10'b1100011000;
mem2[10513] = 10'b1100011000;
mem2[10514] = 10'b1100011000;
mem2[10515] = 10'b1100011000;
mem2[10516] = 10'b1100011000;
mem2[10517] = 10'b1100011000;
mem2[10518] = 10'b1100011000;
mem2[10519] = 10'b1100011000;
mem2[10520] = 10'b1100011001;
mem2[10521] = 10'b1100011001;
mem2[10522] = 10'b1100011001;
mem2[10523] = 10'b1100011001;
mem2[10524] = 10'b1100011001;
mem2[10525] = 10'b1100011001;
mem2[10526] = 10'b1100011001;
mem2[10527] = 10'b1100011001;
mem2[10528] = 10'b1100011001;
mem2[10529] = 10'b1100011001;
mem2[10530] = 10'b1100011001;
mem2[10531] = 10'b1100011001;
mem2[10532] = 10'b1100011010;
mem2[10533] = 10'b1100011010;
mem2[10534] = 10'b1100011010;
mem2[10535] = 10'b1100011010;
mem2[10536] = 10'b1100011010;
mem2[10537] = 10'b1100011010;
mem2[10538] = 10'b1100011010;
mem2[10539] = 10'b1100011010;
mem2[10540] = 10'b1100011010;
mem2[10541] = 10'b1100011010;
mem2[10542] = 10'b1100011010;
mem2[10543] = 10'b1100011011;
mem2[10544] = 10'b1100011011;
mem2[10545] = 10'b1100011011;
mem2[10546] = 10'b1100011011;
mem2[10547] = 10'b1100011011;
mem2[10548] = 10'b1100011011;
mem2[10549] = 10'b1100011011;
mem2[10550] = 10'b1100011011;
mem2[10551] = 10'b1100011011;
mem2[10552] = 10'b1100011011;
mem2[10553] = 10'b1100011011;
mem2[10554] = 10'b1100011011;
mem2[10555] = 10'b1100011100;
mem2[10556] = 10'b1100011100;
mem2[10557] = 10'b1100011100;
mem2[10558] = 10'b1100011100;
mem2[10559] = 10'b1100011100;
mem2[10560] = 10'b1100011100;
mem2[10561] = 10'b1100011100;
mem2[10562] = 10'b1100011100;
mem2[10563] = 10'b1100011100;
mem2[10564] = 10'b1100011100;
mem2[10565] = 10'b1100011100;
mem2[10566] = 10'b1100011101;
mem2[10567] = 10'b1100011101;
mem2[10568] = 10'b1100011101;
mem2[10569] = 10'b1100011101;
mem2[10570] = 10'b1100011101;
mem2[10571] = 10'b1100011101;
mem2[10572] = 10'b1100011101;
mem2[10573] = 10'b1100011101;
mem2[10574] = 10'b1100011101;
mem2[10575] = 10'b1100011101;
mem2[10576] = 10'b1100011101;
mem2[10577] = 10'b1100011101;
mem2[10578] = 10'b1100011110;
mem2[10579] = 10'b1100011110;
mem2[10580] = 10'b1100011110;
mem2[10581] = 10'b1100011110;
mem2[10582] = 10'b1100011110;
mem2[10583] = 10'b1100011110;
mem2[10584] = 10'b1100011110;
mem2[10585] = 10'b1100011110;
mem2[10586] = 10'b1100011110;
mem2[10587] = 10'b1100011110;
mem2[10588] = 10'b1100011110;
mem2[10589] = 10'b1100011111;
mem2[10590] = 10'b1100011111;
mem2[10591] = 10'b1100011111;
mem2[10592] = 10'b1100011111;
mem2[10593] = 10'b1100011111;
mem2[10594] = 10'b1100011111;
mem2[10595] = 10'b1100011111;
mem2[10596] = 10'b1100011111;
mem2[10597] = 10'b1100011111;
mem2[10598] = 10'b1100011111;
mem2[10599] = 10'b1100011111;
mem2[10600] = 10'b1100011111;
mem2[10601] = 10'b1100100000;
mem2[10602] = 10'b1100100000;
mem2[10603] = 10'b1100100000;
mem2[10604] = 10'b1100100000;
mem2[10605] = 10'b1100100000;
mem2[10606] = 10'b1100100000;
mem2[10607] = 10'b1100100000;
mem2[10608] = 10'b1100100000;
mem2[10609] = 10'b1100100000;
mem2[10610] = 10'b1100100000;
mem2[10611] = 10'b1100100000;
mem2[10612] = 10'b1100100001;
mem2[10613] = 10'b1100100001;
mem2[10614] = 10'b1100100001;
mem2[10615] = 10'b1100100001;
mem2[10616] = 10'b1100100001;
mem2[10617] = 10'b1100100001;
mem2[10618] = 10'b1100100001;
mem2[10619] = 10'b1100100001;
mem2[10620] = 10'b1100100001;
mem2[10621] = 10'b1100100001;
mem2[10622] = 10'b1100100001;
mem2[10623] = 10'b1100100001;
mem2[10624] = 10'b1100100010;
mem2[10625] = 10'b1100100010;
mem2[10626] = 10'b1100100010;
mem2[10627] = 10'b1100100010;
mem2[10628] = 10'b1100100010;
mem2[10629] = 10'b1100100010;
mem2[10630] = 10'b1100100010;
mem2[10631] = 10'b1100100010;
mem2[10632] = 10'b1100100010;
mem2[10633] = 10'b1100100010;
mem2[10634] = 10'b1100100010;
mem2[10635] = 10'b1100100010;
mem2[10636] = 10'b1100100011;
mem2[10637] = 10'b1100100011;
mem2[10638] = 10'b1100100011;
mem2[10639] = 10'b1100100011;
mem2[10640] = 10'b1100100011;
mem2[10641] = 10'b1100100011;
mem2[10642] = 10'b1100100011;
mem2[10643] = 10'b1100100011;
mem2[10644] = 10'b1100100011;
mem2[10645] = 10'b1100100011;
mem2[10646] = 10'b1100100011;
mem2[10647] = 10'b1100100100;
mem2[10648] = 10'b1100100100;
mem2[10649] = 10'b1100100100;
mem2[10650] = 10'b1100100100;
mem2[10651] = 10'b1100100100;
mem2[10652] = 10'b1100100100;
mem2[10653] = 10'b1100100100;
mem2[10654] = 10'b1100100100;
mem2[10655] = 10'b1100100100;
mem2[10656] = 10'b1100100100;
mem2[10657] = 10'b1100100100;
mem2[10658] = 10'b1100100100;
mem2[10659] = 10'b1100100101;
mem2[10660] = 10'b1100100101;
mem2[10661] = 10'b1100100101;
mem2[10662] = 10'b1100100101;
mem2[10663] = 10'b1100100101;
mem2[10664] = 10'b1100100101;
mem2[10665] = 10'b1100100101;
mem2[10666] = 10'b1100100101;
mem2[10667] = 10'b1100100101;
mem2[10668] = 10'b1100100101;
mem2[10669] = 10'b1100100101;
mem2[10670] = 10'b1100100110;
mem2[10671] = 10'b1100100110;
mem2[10672] = 10'b1100100110;
mem2[10673] = 10'b1100100110;
mem2[10674] = 10'b1100100110;
mem2[10675] = 10'b1100100110;
mem2[10676] = 10'b1100100110;
mem2[10677] = 10'b1100100110;
mem2[10678] = 10'b1100100110;
mem2[10679] = 10'b1100100110;
mem2[10680] = 10'b1100100110;
mem2[10681] = 10'b1100100110;
mem2[10682] = 10'b1100100111;
mem2[10683] = 10'b1100100111;
mem2[10684] = 10'b1100100111;
mem2[10685] = 10'b1100100111;
mem2[10686] = 10'b1100100111;
mem2[10687] = 10'b1100100111;
mem2[10688] = 10'b1100100111;
mem2[10689] = 10'b1100100111;
mem2[10690] = 10'b1100100111;
mem2[10691] = 10'b1100100111;
mem2[10692] = 10'b1100100111;
mem2[10693] = 10'b1100100111;
mem2[10694] = 10'b1100101000;
mem2[10695] = 10'b1100101000;
mem2[10696] = 10'b1100101000;
mem2[10697] = 10'b1100101000;
mem2[10698] = 10'b1100101000;
mem2[10699] = 10'b1100101000;
mem2[10700] = 10'b1100101000;
mem2[10701] = 10'b1100101000;
mem2[10702] = 10'b1100101000;
mem2[10703] = 10'b1100101000;
mem2[10704] = 10'b1100101000;
mem2[10705] = 10'b1100101001;
mem2[10706] = 10'b1100101001;
mem2[10707] = 10'b1100101001;
mem2[10708] = 10'b1100101001;
mem2[10709] = 10'b1100101001;
mem2[10710] = 10'b1100101001;
mem2[10711] = 10'b1100101001;
mem2[10712] = 10'b1100101001;
mem2[10713] = 10'b1100101001;
mem2[10714] = 10'b1100101001;
mem2[10715] = 10'b1100101001;
mem2[10716] = 10'b1100101001;
mem2[10717] = 10'b1100101010;
mem2[10718] = 10'b1100101010;
mem2[10719] = 10'b1100101010;
mem2[10720] = 10'b1100101010;
mem2[10721] = 10'b1100101010;
mem2[10722] = 10'b1100101010;
mem2[10723] = 10'b1100101010;
mem2[10724] = 10'b1100101010;
mem2[10725] = 10'b1100101010;
mem2[10726] = 10'b1100101010;
mem2[10727] = 10'b1100101010;
mem2[10728] = 10'b1100101010;
mem2[10729] = 10'b1100101011;
mem2[10730] = 10'b1100101011;
mem2[10731] = 10'b1100101011;
mem2[10732] = 10'b1100101011;
mem2[10733] = 10'b1100101011;
mem2[10734] = 10'b1100101011;
mem2[10735] = 10'b1100101011;
mem2[10736] = 10'b1100101011;
mem2[10737] = 10'b1100101011;
mem2[10738] = 10'b1100101011;
mem2[10739] = 10'b1100101011;
mem2[10740] = 10'b1100101011;
mem2[10741] = 10'b1100101100;
mem2[10742] = 10'b1100101100;
mem2[10743] = 10'b1100101100;
mem2[10744] = 10'b1100101100;
mem2[10745] = 10'b1100101100;
mem2[10746] = 10'b1100101100;
mem2[10747] = 10'b1100101100;
mem2[10748] = 10'b1100101100;
mem2[10749] = 10'b1100101100;
mem2[10750] = 10'b1100101100;
mem2[10751] = 10'b1100101100;
mem2[10752] = 10'b1100101100;
mem2[10753] = 10'b1100101101;
mem2[10754] = 10'b1100101101;
mem2[10755] = 10'b1100101101;
mem2[10756] = 10'b1100101101;
mem2[10757] = 10'b1100101101;
mem2[10758] = 10'b1100101101;
mem2[10759] = 10'b1100101101;
mem2[10760] = 10'b1100101101;
mem2[10761] = 10'b1100101101;
mem2[10762] = 10'b1100101101;
mem2[10763] = 10'b1100101101;
mem2[10764] = 10'b1100101110;
mem2[10765] = 10'b1100101110;
mem2[10766] = 10'b1100101110;
mem2[10767] = 10'b1100101110;
mem2[10768] = 10'b1100101110;
mem2[10769] = 10'b1100101110;
mem2[10770] = 10'b1100101110;
mem2[10771] = 10'b1100101110;
mem2[10772] = 10'b1100101110;
mem2[10773] = 10'b1100101110;
mem2[10774] = 10'b1100101110;
mem2[10775] = 10'b1100101110;
mem2[10776] = 10'b1100101111;
mem2[10777] = 10'b1100101111;
mem2[10778] = 10'b1100101111;
mem2[10779] = 10'b1100101111;
mem2[10780] = 10'b1100101111;
mem2[10781] = 10'b1100101111;
mem2[10782] = 10'b1100101111;
mem2[10783] = 10'b1100101111;
mem2[10784] = 10'b1100101111;
mem2[10785] = 10'b1100101111;
mem2[10786] = 10'b1100101111;
mem2[10787] = 10'b1100101111;
mem2[10788] = 10'b1100110000;
mem2[10789] = 10'b1100110000;
mem2[10790] = 10'b1100110000;
mem2[10791] = 10'b1100110000;
mem2[10792] = 10'b1100110000;
mem2[10793] = 10'b1100110000;
mem2[10794] = 10'b1100110000;
mem2[10795] = 10'b1100110000;
mem2[10796] = 10'b1100110000;
mem2[10797] = 10'b1100110000;
mem2[10798] = 10'b1100110000;
mem2[10799] = 10'b1100110000;
mem2[10800] = 10'b1100110001;
mem2[10801] = 10'b1100110001;
mem2[10802] = 10'b1100110001;
mem2[10803] = 10'b1100110001;
mem2[10804] = 10'b1100110001;
mem2[10805] = 10'b1100110001;
mem2[10806] = 10'b1100110001;
mem2[10807] = 10'b1100110001;
mem2[10808] = 10'b1100110001;
mem2[10809] = 10'b1100110001;
mem2[10810] = 10'b1100110001;
mem2[10811] = 10'b1100110001;
mem2[10812] = 10'b1100110010;
mem2[10813] = 10'b1100110010;
mem2[10814] = 10'b1100110010;
mem2[10815] = 10'b1100110010;
mem2[10816] = 10'b1100110010;
mem2[10817] = 10'b1100110010;
mem2[10818] = 10'b1100110010;
mem2[10819] = 10'b1100110010;
mem2[10820] = 10'b1100110010;
mem2[10821] = 10'b1100110010;
mem2[10822] = 10'b1100110010;
mem2[10823] = 10'b1100110010;
mem2[10824] = 10'b1100110011;
mem2[10825] = 10'b1100110011;
mem2[10826] = 10'b1100110011;
mem2[10827] = 10'b1100110011;
mem2[10828] = 10'b1100110011;
mem2[10829] = 10'b1100110011;
mem2[10830] = 10'b1100110011;
mem2[10831] = 10'b1100110011;
mem2[10832] = 10'b1100110011;
mem2[10833] = 10'b1100110011;
mem2[10834] = 10'b1100110011;
mem2[10835] = 10'b1100110011;
mem2[10836] = 10'b1100110100;
mem2[10837] = 10'b1100110100;
mem2[10838] = 10'b1100110100;
mem2[10839] = 10'b1100110100;
mem2[10840] = 10'b1100110100;
mem2[10841] = 10'b1100110100;
mem2[10842] = 10'b1100110100;
mem2[10843] = 10'b1100110100;
mem2[10844] = 10'b1100110100;
mem2[10845] = 10'b1100110100;
mem2[10846] = 10'b1100110100;
mem2[10847] = 10'b1100110100;
mem2[10848] = 10'b1100110101;
mem2[10849] = 10'b1100110101;
mem2[10850] = 10'b1100110101;
mem2[10851] = 10'b1100110101;
mem2[10852] = 10'b1100110101;
mem2[10853] = 10'b1100110101;
mem2[10854] = 10'b1100110101;
mem2[10855] = 10'b1100110101;
mem2[10856] = 10'b1100110101;
mem2[10857] = 10'b1100110101;
mem2[10858] = 10'b1100110101;
mem2[10859] = 10'b1100110101;
mem2[10860] = 10'b1100110110;
mem2[10861] = 10'b1100110110;
mem2[10862] = 10'b1100110110;
mem2[10863] = 10'b1100110110;
mem2[10864] = 10'b1100110110;
mem2[10865] = 10'b1100110110;
mem2[10866] = 10'b1100110110;
mem2[10867] = 10'b1100110110;
mem2[10868] = 10'b1100110110;
mem2[10869] = 10'b1100110110;
mem2[10870] = 10'b1100110110;
mem2[10871] = 10'b1100110110;
mem2[10872] = 10'b1100110111;
mem2[10873] = 10'b1100110111;
mem2[10874] = 10'b1100110111;
mem2[10875] = 10'b1100110111;
mem2[10876] = 10'b1100110111;
mem2[10877] = 10'b1100110111;
mem2[10878] = 10'b1100110111;
mem2[10879] = 10'b1100110111;
mem2[10880] = 10'b1100110111;
mem2[10881] = 10'b1100110111;
mem2[10882] = 10'b1100110111;
mem2[10883] = 10'b1100110111;
mem2[10884] = 10'b1100111000;
mem2[10885] = 10'b1100111000;
mem2[10886] = 10'b1100111000;
mem2[10887] = 10'b1100111000;
mem2[10888] = 10'b1100111000;
mem2[10889] = 10'b1100111000;
mem2[10890] = 10'b1100111000;
mem2[10891] = 10'b1100111000;
mem2[10892] = 10'b1100111000;
mem2[10893] = 10'b1100111000;
mem2[10894] = 10'b1100111000;
mem2[10895] = 10'b1100111000;
mem2[10896] = 10'b1100111001;
mem2[10897] = 10'b1100111001;
mem2[10898] = 10'b1100111001;
mem2[10899] = 10'b1100111001;
mem2[10900] = 10'b1100111001;
mem2[10901] = 10'b1100111001;
mem2[10902] = 10'b1100111001;
mem2[10903] = 10'b1100111001;
mem2[10904] = 10'b1100111001;
mem2[10905] = 10'b1100111001;
mem2[10906] = 10'b1100111001;
mem2[10907] = 10'b1100111001;
mem2[10908] = 10'b1100111010;
mem2[10909] = 10'b1100111010;
mem2[10910] = 10'b1100111010;
mem2[10911] = 10'b1100111010;
mem2[10912] = 10'b1100111010;
mem2[10913] = 10'b1100111010;
mem2[10914] = 10'b1100111010;
mem2[10915] = 10'b1100111010;
mem2[10916] = 10'b1100111010;
mem2[10917] = 10'b1100111010;
mem2[10918] = 10'b1100111010;
mem2[10919] = 10'b1100111010;
mem2[10920] = 10'b1100111011;
mem2[10921] = 10'b1100111011;
mem2[10922] = 10'b1100111011;
mem2[10923] = 10'b1100111011;
mem2[10924] = 10'b1100111011;
mem2[10925] = 10'b1100111011;
mem2[10926] = 10'b1100111011;
mem2[10927] = 10'b1100111011;
mem2[10928] = 10'b1100111011;
mem2[10929] = 10'b1100111011;
mem2[10930] = 10'b1100111011;
mem2[10931] = 10'b1100111011;
mem2[10932] = 10'b1100111100;
mem2[10933] = 10'b1100111100;
mem2[10934] = 10'b1100111100;
mem2[10935] = 10'b1100111100;
mem2[10936] = 10'b1100111100;
mem2[10937] = 10'b1100111100;
mem2[10938] = 10'b1100111100;
mem2[10939] = 10'b1100111100;
mem2[10940] = 10'b1100111100;
mem2[10941] = 10'b1100111100;
mem2[10942] = 10'b1100111100;
mem2[10943] = 10'b1100111100;
mem2[10944] = 10'b1100111101;
mem2[10945] = 10'b1100111101;
mem2[10946] = 10'b1100111101;
mem2[10947] = 10'b1100111101;
mem2[10948] = 10'b1100111101;
mem2[10949] = 10'b1100111101;
mem2[10950] = 10'b1100111101;
mem2[10951] = 10'b1100111101;
mem2[10952] = 10'b1100111101;
mem2[10953] = 10'b1100111101;
mem2[10954] = 10'b1100111101;
mem2[10955] = 10'b1100111101;
mem2[10956] = 10'b1100111110;
mem2[10957] = 10'b1100111110;
mem2[10958] = 10'b1100111110;
mem2[10959] = 10'b1100111110;
mem2[10960] = 10'b1100111110;
mem2[10961] = 10'b1100111110;
mem2[10962] = 10'b1100111110;
mem2[10963] = 10'b1100111110;
mem2[10964] = 10'b1100111110;
mem2[10965] = 10'b1100111110;
mem2[10966] = 10'b1100111110;
mem2[10967] = 10'b1100111110;
mem2[10968] = 10'b1100111110;
mem2[10969] = 10'b1100111111;
mem2[10970] = 10'b1100111111;
mem2[10971] = 10'b1100111111;
mem2[10972] = 10'b1100111111;
mem2[10973] = 10'b1100111111;
mem2[10974] = 10'b1100111111;
mem2[10975] = 10'b1100111111;
mem2[10976] = 10'b1100111111;
mem2[10977] = 10'b1100111111;
mem2[10978] = 10'b1100111111;
mem2[10979] = 10'b1100111111;
mem2[10980] = 10'b1100111111;
mem2[10981] = 10'b1101000000;
mem2[10982] = 10'b1101000000;
mem2[10983] = 10'b1101000000;
mem2[10984] = 10'b1101000000;
mem2[10985] = 10'b1101000000;
mem2[10986] = 10'b1101000000;
mem2[10987] = 10'b1101000000;
mem2[10988] = 10'b1101000000;
mem2[10989] = 10'b1101000000;
mem2[10990] = 10'b1101000000;
mem2[10991] = 10'b1101000000;
mem2[10992] = 10'b1101000000;
mem2[10993] = 10'b1101000001;
mem2[10994] = 10'b1101000001;
mem2[10995] = 10'b1101000001;
mem2[10996] = 10'b1101000001;
mem2[10997] = 10'b1101000001;
mem2[10998] = 10'b1101000001;
mem2[10999] = 10'b1101000001;
mem2[11000] = 10'b1101000001;
mem2[11001] = 10'b1101000001;
mem2[11002] = 10'b1101000001;
mem2[11003] = 10'b1101000001;
mem2[11004] = 10'b1101000001;
mem2[11005] = 10'b1101000010;
mem2[11006] = 10'b1101000010;
mem2[11007] = 10'b1101000010;
mem2[11008] = 10'b1101000010;
mem2[11009] = 10'b1101000010;
mem2[11010] = 10'b1101000010;
mem2[11011] = 10'b1101000010;
mem2[11012] = 10'b1101000010;
mem2[11013] = 10'b1101000010;
mem2[11014] = 10'b1101000010;
mem2[11015] = 10'b1101000010;
mem2[11016] = 10'b1101000010;
mem2[11017] = 10'b1101000010;
mem2[11018] = 10'b1101000011;
mem2[11019] = 10'b1101000011;
mem2[11020] = 10'b1101000011;
mem2[11021] = 10'b1101000011;
mem2[11022] = 10'b1101000011;
mem2[11023] = 10'b1101000011;
mem2[11024] = 10'b1101000011;
mem2[11025] = 10'b1101000011;
mem2[11026] = 10'b1101000011;
mem2[11027] = 10'b1101000011;
mem2[11028] = 10'b1101000011;
mem2[11029] = 10'b1101000011;
mem2[11030] = 10'b1101000100;
mem2[11031] = 10'b1101000100;
mem2[11032] = 10'b1101000100;
mem2[11033] = 10'b1101000100;
mem2[11034] = 10'b1101000100;
mem2[11035] = 10'b1101000100;
mem2[11036] = 10'b1101000100;
mem2[11037] = 10'b1101000100;
mem2[11038] = 10'b1101000100;
mem2[11039] = 10'b1101000100;
mem2[11040] = 10'b1101000100;
mem2[11041] = 10'b1101000100;
mem2[11042] = 10'b1101000101;
mem2[11043] = 10'b1101000101;
mem2[11044] = 10'b1101000101;
mem2[11045] = 10'b1101000101;
mem2[11046] = 10'b1101000101;
mem2[11047] = 10'b1101000101;
mem2[11048] = 10'b1101000101;
mem2[11049] = 10'b1101000101;
mem2[11050] = 10'b1101000101;
mem2[11051] = 10'b1101000101;
mem2[11052] = 10'b1101000101;
mem2[11053] = 10'b1101000101;
mem2[11054] = 10'b1101000101;
mem2[11055] = 10'b1101000110;
mem2[11056] = 10'b1101000110;
mem2[11057] = 10'b1101000110;
mem2[11058] = 10'b1101000110;
mem2[11059] = 10'b1101000110;
mem2[11060] = 10'b1101000110;
mem2[11061] = 10'b1101000110;
mem2[11062] = 10'b1101000110;
mem2[11063] = 10'b1101000110;
mem2[11064] = 10'b1101000110;
mem2[11065] = 10'b1101000110;
mem2[11066] = 10'b1101000110;
mem2[11067] = 10'b1101000111;
mem2[11068] = 10'b1101000111;
mem2[11069] = 10'b1101000111;
mem2[11070] = 10'b1101000111;
mem2[11071] = 10'b1101000111;
mem2[11072] = 10'b1101000111;
mem2[11073] = 10'b1101000111;
mem2[11074] = 10'b1101000111;
mem2[11075] = 10'b1101000111;
mem2[11076] = 10'b1101000111;
mem2[11077] = 10'b1101000111;
mem2[11078] = 10'b1101000111;
mem2[11079] = 10'b1101001000;
mem2[11080] = 10'b1101001000;
mem2[11081] = 10'b1101001000;
mem2[11082] = 10'b1101001000;
mem2[11083] = 10'b1101001000;
mem2[11084] = 10'b1101001000;
mem2[11085] = 10'b1101001000;
mem2[11086] = 10'b1101001000;
mem2[11087] = 10'b1101001000;
mem2[11088] = 10'b1101001000;
mem2[11089] = 10'b1101001000;
mem2[11090] = 10'b1101001000;
mem2[11091] = 10'b1101001000;
mem2[11092] = 10'b1101001001;
mem2[11093] = 10'b1101001001;
mem2[11094] = 10'b1101001001;
mem2[11095] = 10'b1101001001;
mem2[11096] = 10'b1101001001;
mem2[11097] = 10'b1101001001;
mem2[11098] = 10'b1101001001;
mem2[11099] = 10'b1101001001;
mem2[11100] = 10'b1101001001;
mem2[11101] = 10'b1101001001;
mem2[11102] = 10'b1101001001;
mem2[11103] = 10'b1101001001;
mem2[11104] = 10'b1101001010;
mem2[11105] = 10'b1101001010;
mem2[11106] = 10'b1101001010;
mem2[11107] = 10'b1101001010;
mem2[11108] = 10'b1101001010;
mem2[11109] = 10'b1101001010;
mem2[11110] = 10'b1101001010;
mem2[11111] = 10'b1101001010;
mem2[11112] = 10'b1101001010;
mem2[11113] = 10'b1101001010;
mem2[11114] = 10'b1101001010;
mem2[11115] = 10'b1101001010;
mem2[11116] = 10'b1101001010;
mem2[11117] = 10'b1101001011;
mem2[11118] = 10'b1101001011;
mem2[11119] = 10'b1101001011;
mem2[11120] = 10'b1101001011;
mem2[11121] = 10'b1101001011;
mem2[11122] = 10'b1101001011;
mem2[11123] = 10'b1101001011;
mem2[11124] = 10'b1101001011;
mem2[11125] = 10'b1101001011;
mem2[11126] = 10'b1101001011;
mem2[11127] = 10'b1101001011;
mem2[11128] = 10'b1101001011;
mem2[11129] = 10'b1101001100;
mem2[11130] = 10'b1101001100;
mem2[11131] = 10'b1101001100;
mem2[11132] = 10'b1101001100;
mem2[11133] = 10'b1101001100;
mem2[11134] = 10'b1101001100;
mem2[11135] = 10'b1101001100;
mem2[11136] = 10'b1101001100;
mem2[11137] = 10'b1101001100;
mem2[11138] = 10'b1101001100;
mem2[11139] = 10'b1101001100;
mem2[11140] = 10'b1101001100;
mem2[11141] = 10'b1101001100;
mem2[11142] = 10'b1101001101;
mem2[11143] = 10'b1101001101;
mem2[11144] = 10'b1101001101;
mem2[11145] = 10'b1101001101;
mem2[11146] = 10'b1101001101;
mem2[11147] = 10'b1101001101;
mem2[11148] = 10'b1101001101;
mem2[11149] = 10'b1101001101;
mem2[11150] = 10'b1101001101;
mem2[11151] = 10'b1101001101;
mem2[11152] = 10'b1101001101;
mem2[11153] = 10'b1101001101;
mem2[11154] = 10'b1101001101;
mem2[11155] = 10'b1101001110;
mem2[11156] = 10'b1101001110;
mem2[11157] = 10'b1101001110;
mem2[11158] = 10'b1101001110;
mem2[11159] = 10'b1101001110;
mem2[11160] = 10'b1101001110;
mem2[11161] = 10'b1101001110;
mem2[11162] = 10'b1101001110;
mem2[11163] = 10'b1101001110;
mem2[11164] = 10'b1101001110;
mem2[11165] = 10'b1101001110;
mem2[11166] = 10'b1101001110;
mem2[11167] = 10'b1101001111;
mem2[11168] = 10'b1101001111;
mem2[11169] = 10'b1101001111;
mem2[11170] = 10'b1101001111;
mem2[11171] = 10'b1101001111;
mem2[11172] = 10'b1101001111;
mem2[11173] = 10'b1101001111;
mem2[11174] = 10'b1101001111;
mem2[11175] = 10'b1101001111;
mem2[11176] = 10'b1101001111;
mem2[11177] = 10'b1101001111;
mem2[11178] = 10'b1101001111;
mem2[11179] = 10'b1101001111;
mem2[11180] = 10'b1101010000;
mem2[11181] = 10'b1101010000;
mem2[11182] = 10'b1101010000;
mem2[11183] = 10'b1101010000;
mem2[11184] = 10'b1101010000;
mem2[11185] = 10'b1101010000;
mem2[11186] = 10'b1101010000;
mem2[11187] = 10'b1101010000;
mem2[11188] = 10'b1101010000;
mem2[11189] = 10'b1101010000;
mem2[11190] = 10'b1101010000;
mem2[11191] = 10'b1101010000;
mem2[11192] = 10'b1101010001;
mem2[11193] = 10'b1101010001;
mem2[11194] = 10'b1101010001;
mem2[11195] = 10'b1101010001;
mem2[11196] = 10'b1101010001;
mem2[11197] = 10'b1101010001;
mem2[11198] = 10'b1101010001;
mem2[11199] = 10'b1101010001;
mem2[11200] = 10'b1101010001;
mem2[11201] = 10'b1101010001;
mem2[11202] = 10'b1101010001;
mem2[11203] = 10'b1101010001;
mem2[11204] = 10'b1101010001;
mem2[11205] = 10'b1101010010;
mem2[11206] = 10'b1101010010;
mem2[11207] = 10'b1101010010;
mem2[11208] = 10'b1101010010;
mem2[11209] = 10'b1101010010;
mem2[11210] = 10'b1101010010;
mem2[11211] = 10'b1101010010;
mem2[11212] = 10'b1101010010;
mem2[11213] = 10'b1101010010;
mem2[11214] = 10'b1101010010;
mem2[11215] = 10'b1101010010;
mem2[11216] = 10'b1101010010;
mem2[11217] = 10'b1101010010;
mem2[11218] = 10'b1101010011;
mem2[11219] = 10'b1101010011;
mem2[11220] = 10'b1101010011;
mem2[11221] = 10'b1101010011;
mem2[11222] = 10'b1101010011;
mem2[11223] = 10'b1101010011;
mem2[11224] = 10'b1101010011;
mem2[11225] = 10'b1101010011;
mem2[11226] = 10'b1101010011;
mem2[11227] = 10'b1101010011;
mem2[11228] = 10'b1101010011;
mem2[11229] = 10'b1101010011;
mem2[11230] = 10'b1101010011;
mem2[11231] = 10'b1101010100;
mem2[11232] = 10'b1101010100;
mem2[11233] = 10'b1101010100;
mem2[11234] = 10'b1101010100;
mem2[11235] = 10'b1101010100;
mem2[11236] = 10'b1101010100;
mem2[11237] = 10'b1101010100;
mem2[11238] = 10'b1101010100;
mem2[11239] = 10'b1101010100;
mem2[11240] = 10'b1101010100;
mem2[11241] = 10'b1101010100;
mem2[11242] = 10'b1101010100;
mem2[11243] = 10'b1101010101;
mem2[11244] = 10'b1101010101;
mem2[11245] = 10'b1101010101;
mem2[11246] = 10'b1101010101;
mem2[11247] = 10'b1101010101;
mem2[11248] = 10'b1101010101;
mem2[11249] = 10'b1101010101;
mem2[11250] = 10'b1101010101;
mem2[11251] = 10'b1101010101;
mem2[11252] = 10'b1101010101;
mem2[11253] = 10'b1101010101;
mem2[11254] = 10'b1101010101;
mem2[11255] = 10'b1101010101;
mem2[11256] = 10'b1101010110;
mem2[11257] = 10'b1101010110;
mem2[11258] = 10'b1101010110;
mem2[11259] = 10'b1101010110;
mem2[11260] = 10'b1101010110;
mem2[11261] = 10'b1101010110;
mem2[11262] = 10'b1101010110;
mem2[11263] = 10'b1101010110;
mem2[11264] = 10'b1101010110;
mem2[11265] = 10'b1101010110;
mem2[11266] = 10'b1101010110;
mem2[11267] = 10'b1101010110;
mem2[11268] = 10'b1101010110;
mem2[11269] = 10'b1101010111;
mem2[11270] = 10'b1101010111;
mem2[11271] = 10'b1101010111;
mem2[11272] = 10'b1101010111;
mem2[11273] = 10'b1101010111;
mem2[11274] = 10'b1101010111;
mem2[11275] = 10'b1101010111;
mem2[11276] = 10'b1101010111;
mem2[11277] = 10'b1101010111;
mem2[11278] = 10'b1101010111;
mem2[11279] = 10'b1101010111;
mem2[11280] = 10'b1101010111;
mem2[11281] = 10'b1101010111;
mem2[11282] = 10'b1101011000;
mem2[11283] = 10'b1101011000;
mem2[11284] = 10'b1101011000;
mem2[11285] = 10'b1101011000;
mem2[11286] = 10'b1101011000;
mem2[11287] = 10'b1101011000;
mem2[11288] = 10'b1101011000;
mem2[11289] = 10'b1101011000;
mem2[11290] = 10'b1101011000;
mem2[11291] = 10'b1101011000;
mem2[11292] = 10'b1101011000;
mem2[11293] = 10'b1101011000;
mem2[11294] = 10'b1101011000;
mem2[11295] = 10'b1101011001;
mem2[11296] = 10'b1101011001;
mem2[11297] = 10'b1101011001;
mem2[11298] = 10'b1101011001;
mem2[11299] = 10'b1101011001;
mem2[11300] = 10'b1101011001;
mem2[11301] = 10'b1101011001;
mem2[11302] = 10'b1101011001;
mem2[11303] = 10'b1101011001;
mem2[11304] = 10'b1101011001;
mem2[11305] = 10'b1101011001;
mem2[11306] = 10'b1101011001;
mem2[11307] = 10'b1101011001;
mem2[11308] = 10'b1101011010;
mem2[11309] = 10'b1101011010;
mem2[11310] = 10'b1101011010;
mem2[11311] = 10'b1101011010;
mem2[11312] = 10'b1101011010;
mem2[11313] = 10'b1101011010;
mem2[11314] = 10'b1101011010;
mem2[11315] = 10'b1101011010;
mem2[11316] = 10'b1101011010;
mem2[11317] = 10'b1101011010;
mem2[11318] = 10'b1101011010;
mem2[11319] = 10'b1101011010;
mem2[11320] = 10'b1101011010;
mem2[11321] = 10'b1101011011;
mem2[11322] = 10'b1101011011;
mem2[11323] = 10'b1101011011;
mem2[11324] = 10'b1101011011;
mem2[11325] = 10'b1101011011;
mem2[11326] = 10'b1101011011;
mem2[11327] = 10'b1101011011;
mem2[11328] = 10'b1101011011;
mem2[11329] = 10'b1101011011;
mem2[11330] = 10'b1101011011;
mem2[11331] = 10'b1101011011;
mem2[11332] = 10'b1101011011;
mem2[11333] = 10'b1101011011;
mem2[11334] = 10'b1101011100;
mem2[11335] = 10'b1101011100;
mem2[11336] = 10'b1101011100;
mem2[11337] = 10'b1101011100;
mem2[11338] = 10'b1101011100;
mem2[11339] = 10'b1101011100;
mem2[11340] = 10'b1101011100;
mem2[11341] = 10'b1101011100;
mem2[11342] = 10'b1101011100;
mem2[11343] = 10'b1101011100;
mem2[11344] = 10'b1101011100;
mem2[11345] = 10'b1101011100;
mem2[11346] = 10'b1101011100;
mem2[11347] = 10'b1101011101;
mem2[11348] = 10'b1101011101;
mem2[11349] = 10'b1101011101;
mem2[11350] = 10'b1101011101;
mem2[11351] = 10'b1101011101;
mem2[11352] = 10'b1101011101;
mem2[11353] = 10'b1101011101;
mem2[11354] = 10'b1101011101;
mem2[11355] = 10'b1101011101;
mem2[11356] = 10'b1101011101;
mem2[11357] = 10'b1101011101;
mem2[11358] = 10'b1101011101;
mem2[11359] = 10'b1101011101;
mem2[11360] = 10'b1101011110;
mem2[11361] = 10'b1101011110;
mem2[11362] = 10'b1101011110;
mem2[11363] = 10'b1101011110;
mem2[11364] = 10'b1101011110;
mem2[11365] = 10'b1101011110;
mem2[11366] = 10'b1101011110;
mem2[11367] = 10'b1101011110;
mem2[11368] = 10'b1101011110;
mem2[11369] = 10'b1101011110;
mem2[11370] = 10'b1101011110;
mem2[11371] = 10'b1101011110;
mem2[11372] = 10'b1101011110;
mem2[11373] = 10'b1101011111;
mem2[11374] = 10'b1101011111;
mem2[11375] = 10'b1101011111;
mem2[11376] = 10'b1101011111;
mem2[11377] = 10'b1101011111;
mem2[11378] = 10'b1101011111;
mem2[11379] = 10'b1101011111;
mem2[11380] = 10'b1101011111;
mem2[11381] = 10'b1101011111;
mem2[11382] = 10'b1101011111;
mem2[11383] = 10'b1101011111;
mem2[11384] = 10'b1101011111;
mem2[11385] = 10'b1101011111;
mem2[11386] = 10'b1101100000;
mem2[11387] = 10'b1101100000;
mem2[11388] = 10'b1101100000;
mem2[11389] = 10'b1101100000;
mem2[11390] = 10'b1101100000;
mem2[11391] = 10'b1101100000;
mem2[11392] = 10'b1101100000;
mem2[11393] = 10'b1101100000;
mem2[11394] = 10'b1101100000;
mem2[11395] = 10'b1101100000;
mem2[11396] = 10'b1101100000;
mem2[11397] = 10'b1101100000;
mem2[11398] = 10'b1101100000;
mem2[11399] = 10'b1101100001;
mem2[11400] = 10'b1101100001;
mem2[11401] = 10'b1101100001;
mem2[11402] = 10'b1101100001;
mem2[11403] = 10'b1101100001;
mem2[11404] = 10'b1101100001;
mem2[11405] = 10'b1101100001;
mem2[11406] = 10'b1101100001;
mem2[11407] = 10'b1101100001;
mem2[11408] = 10'b1101100001;
mem2[11409] = 10'b1101100001;
mem2[11410] = 10'b1101100001;
mem2[11411] = 10'b1101100001;
mem2[11412] = 10'b1101100010;
mem2[11413] = 10'b1101100010;
mem2[11414] = 10'b1101100010;
mem2[11415] = 10'b1101100010;
mem2[11416] = 10'b1101100010;
mem2[11417] = 10'b1101100010;
mem2[11418] = 10'b1101100010;
mem2[11419] = 10'b1101100010;
mem2[11420] = 10'b1101100010;
mem2[11421] = 10'b1101100010;
mem2[11422] = 10'b1101100010;
mem2[11423] = 10'b1101100010;
mem2[11424] = 10'b1101100010;
mem2[11425] = 10'b1101100010;
mem2[11426] = 10'b1101100011;
mem2[11427] = 10'b1101100011;
mem2[11428] = 10'b1101100011;
mem2[11429] = 10'b1101100011;
mem2[11430] = 10'b1101100011;
mem2[11431] = 10'b1101100011;
mem2[11432] = 10'b1101100011;
mem2[11433] = 10'b1101100011;
mem2[11434] = 10'b1101100011;
mem2[11435] = 10'b1101100011;
mem2[11436] = 10'b1101100011;
mem2[11437] = 10'b1101100011;
mem2[11438] = 10'b1101100011;
mem2[11439] = 10'b1101100100;
mem2[11440] = 10'b1101100100;
mem2[11441] = 10'b1101100100;
mem2[11442] = 10'b1101100100;
mem2[11443] = 10'b1101100100;
mem2[11444] = 10'b1101100100;
mem2[11445] = 10'b1101100100;
mem2[11446] = 10'b1101100100;
mem2[11447] = 10'b1101100100;
mem2[11448] = 10'b1101100100;
mem2[11449] = 10'b1101100100;
mem2[11450] = 10'b1101100100;
mem2[11451] = 10'b1101100100;
mem2[11452] = 10'b1101100101;
mem2[11453] = 10'b1101100101;
mem2[11454] = 10'b1101100101;
mem2[11455] = 10'b1101100101;
mem2[11456] = 10'b1101100101;
mem2[11457] = 10'b1101100101;
mem2[11458] = 10'b1101100101;
mem2[11459] = 10'b1101100101;
mem2[11460] = 10'b1101100101;
mem2[11461] = 10'b1101100101;
mem2[11462] = 10'b1101100101;
mem2[11463] = 10'b1101100101;
mem2[11464] = 10'b1101100101;
mem2[11465] = 10'b1101100101;
mem2[11466] = 10'b1101100110;
mem2[11467] = 10'b1101100110;
mem2[11468] = 10'b1101100110;
mem2[11469] = 10'b1101100110;
mem2[11470] = 10'b1101100110;
mem2[11471] = 10'b1101100110;
mem2[11472] = 10'b1101100110;
mem2[11473] = 10'b1101100110;
mem2[11474] = 10'b1101100110;
mem2[11475] = 10'b1101100110;
mem2[11476] = 10'b1101100110;
mem2[11477] = 10'b1101100110;
mem2[11478] = 10'b1101100110;
mem2[11479] = 10'b1101100111;
mem2[11480] = 10'b1101100111;
mem2[11481] = 10'b1101100111;
mem2[11482] = 10'b1101100111;
mem2[11483] = 10'b1101100111;
mem2[11484] = 10'b1101100111;
mem2[11485] = 10'b1101100111;
mem2[11486] = 10'b1101100111;
mem2[11487] = 10'b1101100111;
mem2[11488] = 10'b1101100111;
mem2[11489] = 10'b1101100111;
mem2[11490] = 10'b1101100111;
mem2[11491] = 10'b1101100111;
mem2[11492] = 10'b1101101000;
mem2[11493] = 10'b1101101000;
mem2[11494] = 10'b1101101000;
mem2[11495] = 10'b1101101000;
mem2[11496] = 10'b1101101000;
mem2[11497] = 10'b1101101000;
mem2[11498] = 10'b1101101000;
mem2[11499] = 10'b1101101000;
mem2[11500] = 10'b1101101000;
mem2[11501] = 10'b1101101000;
mem2[11502] = 10'b1101101000;
mem2[11503] = 10'b1101101000;
mem2[11504] = 10'b1101101000;
mem2[11505] = 10'b1101101000;
mem2[11506] = 10'b1101101001;
mem2[11507] = 10'b1101101001;
mem2[11508] = 10'b1101101001;
mem2[11509] = 10'b1101101001;
mem2[11510] = 10'b1101101001;
mem2[11511] = 10'b1101101001;
mem2[11512] = 10'b1101101001;
mem2[11513] = 10'b1101101001;
mem2[11514] = 10'b1101101001;
mem2[11515] = 10'b1101101001;
mem2[11516] = 10'b1101101001;
mem2[11517] = 10'b1101101001;
mem2[11518] = 10'b1101101001;
mem2[11519] = 10'b1101101010;
mem2[11520] = 10'b1101101010;
mem2[11521] = 10'b1101101010;
mem2[11522] = 10'b1101101010;
mem2[11523] = 10'b1101101010;
mem2[11524] = 10'b1101101010;
mem2[11525] = 10'b1101101010;
mem2[11526] = 10'b1101101010;
mem2[11527] = 10'b1101101010;
mem2[11528] = 10'b1101101010;
mem2[11529] = 10'b1101101010;
mem2[11530] = 10'b1101101010;
mem2[11531] = 10'b1101101010;
mem2[11532] = 10'b1101101010;
mem2[11533] = 10'b1101101011;
mem2[11534] = 10'b1101101011;
mem2[11535] = 10'b1101101011;
mem2[11536] = 10'b1101101011;
mem2[11537] = 10'b1101101011;
mem2[11538] = 10'b1101101011;
mem2[11539] = 10'b1101101011;
mem2[11540] = 10'b1101101011;
mem2[11541] = 10'b1101101011;
mem2[11542] = 10'b1101101011;
mem2[11543] = 10'b1101101011;
mem2[11544] = 10'b1101101011;
mem2[11545] = 10'b1101101011;
mem2[11546] = 10'b1101101100;
mem2[11547] = 10'b1101101100;
mem2[11548] = 10'b1101101100;
mem2[11549] = 10'b1101101100;
mem2[11550] = 10'b1101101100;
mem2[11551] = 10'b1101101100;
mem2[11552] = 10'b1101101100;
mem2[11553] = 10'b1101101100;
mem2[11554] = 10'b1101101100;
mem2[11555] = 10'b1101101100;
mem2[11556] = 10'b1101101100;
mem2[11557] = 10'b1101101100;
mem2[11558] = 10'b1101101100;
mem2[11559] = 10'b1101101100;
mem2[11560] = 10'b1101101101;
mem2[11561] = 10'b1101101101;
mem2[11562] = 10'b1101101101;
mem2[11563] = 10'b1101101101;
mem2[11564] = 10'b1101101101;
mem2[11565] = 10'b1101101101;
mem2[11566] = 10'b1101101101;
mem2[11567] = 10'b1101101101;
mem2[11568] = 10'b1101101101;
mem2[11569] = 10'b1101101101;
mem2[11570] = 10'b1101101101;
mem2[11571] = 10'b1101101101;
mem2[11572] = 10'b1101101101;
mem2[11573] = 10'b1101101101;
mem2[11574] = 10'b1101101110;
mem2[11575] = 10'b1101101110;
mem2[11576] = 10'b1101101110;
mem2[11577] = 10'b1101101110;
mem2[11578] = 10'b1101101110;
mem2[11579] = 10'b1101101110;
mem2[11580] = 10'b1101101110;
mem2[11581] = 10'b1101101110;
mem2[11582] = 10'b1101101110;
mem2[11583] = 10'b1101101110;
mem2[11584] = 10'b1101101110;
mem2[11585] = 10'b1101101110;
mem2[11586] = 10'b1101101110;
mem2[11587] = 10'b1101101111;
mem2[11588] = 10'b1101101111;
mem2[11589] = 10'b1101101111;
mem2[11590] = 10'b1101101111;
mem2[11591] = 10'b1101101111;
mem2[11592] = 10'b1101101111;
mem2[11593] = 10'b1101101111;
mem2[11594] = 10'b1101101111;
mem2[11595] = 10'b1101101111;
mem2[11596] = 10'b1101101111;
mem2[11597] = 10'b1101101111;
mem2[11598] = 10'b1101101111;
mem2[11599] = 10'b1101101111;
mem2[11600] = 10'b1101101111;
mem2[11601] = 10'b1101110000;
mem2[11602] = 10'b1101110000;
mem2[11603] = 10'b1101110000;
mem2[11604] = 10'b1101110000;
mem2[11605] = 10'b1101110000;
mem2[11606] = 10'b1101110000;
mem2[11607] = 10'b1101110000;
mem2[11608] = 10'b1101110000;
mem2[11609] = 10'b1101110000;
mem2[11610] = 10'b1101110000;
mem2[11611] = 10'b1101110000;
mem2[11612] = 10'b1101110000;
mem2[11613] = 10'b1101110000;
mem2[11614] = 10'b1101110000;
mem2[11615] = 10'b1101110001;
mem2[11616] = 10'b1101110001;
mem2[11617] = 10'b1101110001;
mem2[11618] = 10'b1101110001;
mem2[11619] = 10'b1101110001;
mem2[11620] = 10'b1101110001;
mem2[11621] = 10'b1101110001;
mem2[11622] = 10'b1101110001;
mem2[11623] = 10'b1101110001;
mem2[11624] = 10'b1101110001;
mem2[11625] = 10'b1101110001;
mem2[11626] = 10'b1101110001;
mem2[11627] = 10'b1101110001;
mem2[11628] = 10'b1101110001;
mem2[11629] = 10'b1101110010;
mem2[11630] = 10'b1101110010;
mem2[11631] = 10'b1101110010;
mem2[11632] = 10'b1101110010;
mem2[11633] = 10'b1101110010;
mem2[11634] = 10'b1101110010;
mem2[11635] = 10'b1101110010;
mem2[11636] = 10'b1101110010;
mem2[11637] = 10'b1101110010;
mem2[11638] = 10'b1101110010;
mem2[11639] = 10'b1101110010;
mem2[11640] = 10'b1101110010;
mem2[11641] = 10'b1101110010;
mem2[11642] = 10'b1101110011;
mem2[11643] = 10'b1101110011;
mem2[11644] = 10'b1101110011;
mem2[11645] = 10'b1101110011;
mem2[11646] = 10'b1101110011;
mem2[11647] = 10'b1101110011;
mem2[11648] = 10'b1101110011;
mem2[11649] = 10'b1101110011;
mem2[11650] = 10'b1101110011;
mem2[11651] = 10'b1101110011;
mem2[11652] = 10'b1101110011;
mem2[11653] = 10'b1101110011;
mem2[11654] = 10'b1101110011;
mem2[11655] = 10'b1101110011;
mem2[11656] = 10'b1101110100;
mem2[11657] = 10'b1101110100;
mem2[11658] = 10'b1101110100;
mem2[11659] = 10'b1101110100;
mem2[11660] = 10'b1101110100;
mem2[11661] = 10'b1101110100;
mem2[11662] = 10'b1101110100;
mem2[11663] = 10'b1101110100;
mem2[11664] = 10'b1101110100;
mem2[11665] = 10'b1101110100;
mem2[11666] = 10'b1101110100;
mem2[11667] = 10'b1101110100;
mem2[11668] = 10'b1101110100;
mem2[11669] = 10'b1101110100;
mem2[11670] = 10'b1101110101;
mem2[11671] = 10'b1101110101;
mem2[11672] = 10'b1101110101;
mem2[11673] = 10'b1101110101;
mem2[11674] = 10'b1101110101;
mem2[11675] = 10'b1101110101;
mem2[11676] = 10'b1101110101;
mem2[11677] = 10'b1101110101;
mem2[11678] = 10'b1101110101;
mem2[11679] = 10'b1101110101;
mem2[11680] = 10'b1101110101;
mem2[11681] = 10'b1101110101;
mem2[11682] = 10'b1101110101;
mem2[11683] = 10'b1101110101;
mem2[11684] = 10'b1101110110;
mem2[11685] = 10'b1101110110;
mem2[11686] = 10'b1101110110;
mem2[11687] = 10'b1101110110;
mem2[11688] = 10'b1101110110;
mem2[11689] = 10'b1101110110;
mem2[11690] = 10'b1101110110;
mem2[11691] = 10'b1101110110;
mem2[11692] = 10'b1101110110;
mem2[11693] = 10'b1101110110;
mem2[11694] = 10'b1101110110;
mem2[11695] = 10'b1101110110;
mem2[11696] = 10'b1101110110;
mem2[11697] = 10'b1101110110;
mem2[11698] = 10'b1101110111;
mem2[11699] = 10'b1101110111;
mem2[11700] = 10'b1101110111;
mem2[11701] = 10'b1101110111;
mem2[11702] = 10'b1101110111;
mem2[11703] = 10'b1101110111;
mem2[11704] = 10'b1101110111;
mem2[11705] = 10'b1101110111;
mem2[11706] = 10'b1101110111;
mem2[11707] = 10'b1101110111;
mem2[11708] = 10'b1101110111;
mem2[11709] = 10'b1101110111;
mem2[11710] = 10'b1101110111;
mem2[11711] = 10'b1101110111;
mem2[11712] = 10'b1101111000;
mem2[11713] = 10'b1101111000;
mem2[11714] = 10'b1101111000;
mem2[11715] = 10'b1101111000;
mem2[11716] = 10'b1101111000;
mem2[11717] = 10'b1101111000;
mem2[11718] = 10'b1101111000;
mem2[11719] = 10'b1101111000;
mem2[11720] = 10'b1101111000;
mem2[11721] = 10'b1101111000;
mem2[11722] = 10'b1101111000;
mem2[11723] = 10'b1101111000;
mem2[11724] = 10'b1101111000;
mem2[11725] = 10'b1101111000;
mem2[11726] = 10'b1101111001;
mem2[11727] = 10'b1101111001;
mem2[11728] = 10'b1101111001;
mem2[11729] = 10'b1101111001;
mem2[11730] = 10'b1101111001;
mem2[11731] = 10'b1101111001;
mem2[11732] = 10'b1101111001;
mem2[11733] = 10'b1101111001;
mem2[11734] = 10'b1101111001;
mem2[11735] = 10'b1101111001;
mem2[11736] = 10'b1101111001;
mem2[11737] = 10'b1101111001;
mem2[11738] = 10'b1101111001;
mem2[11739] = 10'b1101111001;
mem2[11740] = 10'b1101111010;
mem2[11741] = 10'b1101111010;
mem2[11742] = 10'b1101111010;
mem2[11743] = 10'b1101111010;
mem2[11744] = 10'b1101111010;
mem2[11745] = 10'b1101111010;
mem2[11746] = 10'b1101111010;
mem2[11747] = 10'b1101111010;
mem2[11748] = 10'b1101111010;
mem2[11749] = 10'b1101111010;
mem2[11750] = 10'b1101111010;
mem2[11751] = 10'b1101111010;
mem2[11752] = 10'b1101111010;
mem2[11753] = 10'b1101111010;
mem2[11754] = 10'b1101111010;
mem2[11755] = 10'b1101111011;
mem2[11756] = 10'b1101111011;
mem2[11757] = 10'b1101111011;
mem2[11758] = 10'b1101111011;
mem2[11759] = 10'b1101111011;
mem2[11760] = 10'b1101111011;
mem2[11761] = 10'b1101111011;
mem2[11762] = 10'b1101111011;
mem2[11763] = 10'b1101111011;
mem2[11764] = 10'b1101111011;
mem2[11765] = 10'b1101111011;
mem2[11766] = 10'b1101111011;
mem2[11767] = 10'b1101111011;
mem2[11768] = 10'b1101111011;
mem2[11769] = 10'b1101111100;
mem2[11770] = 10'b1101111100;
mem2[11771] = 10'b1101111100;
mem2[11772] = 10'b1101111100;
mem2[11773] = 10'b1101111100;
mem2[11774] = 10'b1101111100;
mem2[11775] = 10'b1101111100;
mem2[11776] = 10'b1101111100;
mem2[11777] = 10'b1101111100;
mem2[11778] = 10'b1101111100;
mem2[11779] = 10'b1101111100;
mem2[11780] = 10'b1101111100;
mem2[11781] = 10'b1101111100;
mem2[11782] = 10'b1101111100;
mem2[11783] = 10'b1101111101;
mem2[11784] = 10'b1101111101;
mem2[11785] = 10'b1101111101;
mem2[11786] = 10'b1101111101;
mem2[11787] = 10'b1101111101;
mem2[11788] = 10'b1101111101;
mem2[11789] = 10'b1101111101;
mem2[11790] = 10'b1101111101;
mem2[11791] = 10'b1101111101;
mem2[11792] = 10'b1101111101;
mem2[11793] = 10'b1101111101;
mem2[11794] = 10'b1101111101;
mem2[11795] = 10'b1101111101;
mem2[11796] = 10'b1101111101;
mem2[11797] = 10'b1101111110;
mem2[11798] = 10'b1101111110;
mem2[11799] = 10'b1101111110;
mem2[11800] = 10'b1101111110;
mem2[11801] = 10'b1101111110;
mem2[11802] = 10'b1101111110;
mem2[11803] = 10'b1101111110;
mem2[11804] = 10'b1101111110;
mem2[11805] = 10'b1101111110;
mem2[11806] = 10'b1101111110;
mem2[11807] = 10'b1101111110;
mem2[11808] = 10'b1101111110;
mem2[11809] = 10'b1101111110;
mem2[11810] = 10'b1101111110;
mem2[11811] = 10'b1101111110;
mem2[11812] = 10'b1101111111;
mem2[11813] = 10'b1101111111;
mem2[11814] = 10'b1101111111;
mem2[11815] = 10'b1101111111;
mem2[11816] = 10'b1101111111;
mem2[11817] = 10'b1101111111;
mem2[11818] = 10'b1101111111;
mem2[11819] = 10'b1101111111;
mem2[11820] = 10'b1101111111;
mem2[11821] = 10'b1101111111;
mem2[11822] = 10'b1101111111;
mem2[11823] = 10'b1101111111;
mem2[11824] = 10'b1101111111;
mem2[11825] = 10'b1101111111;
mem2[11826] = 10'b1110000000;
mem2[11827] = 10'b1110000000;
mem2[11828] = 10'b1110000000;
mem2[11829] = 10'b1110000000;
mem2[11830] = 10'b1110000000;
mem2[11831] = 10'b1110000000;
mem2[11832] = 10'b1110000000;
mem2[11833] = 10'b1110000000;
mem2[11834] = 10'b1110000000;
mem2[11835] = 10'b1110000000;
mem2[11836] = 10'b1110000000;
mem2[11837] = 10'b1110000000;
mem2[11838] = 10'b1110000000;
mem2[11839] = 10'b1110000000;
mem2[11840] = 10'b1110000000;
mem2[11841] = 10'b1110000001;
mem2[11842] = 10'b1110000001;
mem2[11843] = 10'b1110000001;
mem2[11844] = 10'b1110000001;
mem2[11845] = 10'b1110000001;
mem2[11846] = 10'b1110000001;
mem2[11847] = 10'b1110000001;
mem2[11848] = 10'b1110000001;
mem2[11849] = 10'b1110000001;
mem2[11850] = 10'b1110000001;
mem2[11851] = 10'b1110000001;
mem2[11852] = 10'b1110000001;
mem2[11853] = 10'b1110000001;
mem2[11854] = 10'b1110000001;
mem2[11855] = 10'b1110000010;
mem2[11856] = 10'b1110000010;
mem2[11857] = 10'b1110000010;
mem2[11858] = 10'b1110000010;
mem2[11859] = 10'b1110000010;
mem2[11860] = 10'b1110000010;
mem2[11861] = 10'b1110000010;
mem2[11862] = 10'b1110000010;
mem2[11863] = 10'b1110000010;
mem2[11864] = 10'b1110000010;
mem2[11865] = 10'b1110000010;
mem2[11866] = 10'b1110000010;
mem2[11867] = 10'b1110000010;
mem2[11868] = 10'b1110000010;
mem2[11869] = 10'b1110000010;
mem2[11870] = 10'b1110000011;
mem2[11871] = 10'b1110000011;
mem2[11872] = 10'b1110000011;
mem2[11873] = 10'b1110000011;
mem2[11874] = 10'b1110000011;
mem2[11875] = 10'b1110000011;
mem2[11876] = 10'b1110000011;
mem2[11877] = 10'b1110000011;
mem2[11878] = 10'b1110000011;
mem2[11879] = 10'b1110000011;
mem2[11880] = 10'b1110000011;
mem2[11881] = 10'b1110000011;
mem2[11882] = 10'b1110000011;
mem2[11883] = 10'b1110000011;
mem2[11884] = 10'b1110000100;
mem2[11885] = 10'b1110000100;
mem2[11886] = 10'b1110000100;
mem2[11887] = 10'b1110000100;
mem2[11888] = 10'b1110000100;
mem2[11889] = 10'b1110000100;
mem2[11890] = 10'b1110000100;
mem2[11891] = 10'b1110000100;
mem2[11892] = 10'b1110000100;
mem2[11893] = 10'b1110000100;
mem2[11894] = 10'b1110000100;
mem2[11895] = 10'b1110000100;
mem2[11896] = 10'b1110000100;
mem2[11897] = 10'b1110000100;
mem2[11898] = 10'b1110000100;
mem2[11899] = 10'b1110000101;
mem2[11900] = 10'b1110000101;
mem2[11901] = 10'b1110000101;
mem2[11902] = 10'b1110000101;
mem2[11903] = 10'b1110000101;
mem2[11904] = 10'b1110000101;
mem2[11905] = 10'b1110000101;
mem2[11906] = 10'b1110000101;
mem2[11907] = 10'b1110000101;
mem2[11908] = 10'b1110000101;
mem2[11909] = 10'b1110000101;
mem2[11910] = 10'b1110000101;
mem2[11911] = 10'b1110000101;
mem2[11912] = 10'b1110000101;
mem2[11913] = 10'b1110000101;
mem2[11914] = 10'b1110000110;
mem2[11915] = 10'b1110000110;
mem2[11916] = 10'b1110000110;
mem2[11917] = 10'b1110000110;
mem2[11918] = 10'b1110000110;
mem2[11919] = 10'b1110000110;
mem2[11920] = 10'b1110000110;
mem2[11921] = 10'b1110000110;
mem2[11922] = 10'b1110000110;
mem2[11923] = 10'b1110000110;
mem2[11924] = 10'b1110000110;
mem2[11925] = 10'b1110000110;
mem2[11926] = 10'b1110000110;
mem2[11927] = 10'b1110000110;
mem2[11928] = 10'b1110000110;
mem2[11929] = 10'b1110000111;
mem2[11930] = 10'b1110000111;
mem2[11931] = 10'b1110000111;
mem2[11932] = 10'b1110000111;
mem2[11933] = 10'b1110000111;
mem2[11934] = 10'b1110000111;
mem2[11935] = 10'b1110000111;
mem2[11936] = 10'b1110000111;
mem2[11937] = 10'b1110000111;
mem2[11938] = 10'b1110000111;
mem2[11939] = 10'b1110000111;
mem2[11940] = 10'b1110000111;
mem2[11941] = 10'b1110000111;
mem2[11942] = 10'b1110000111;
mem2[11943] = 10'b1110001000;
mem2[11944] = 10'b1110001000;
mem2[11945] = 10'b1110001000;
mem2[11946] = 10'b1110001000;
mem2[11947] = 10'b1110001000;
mem2[11948] = 10'b1110001000;
mem2[11949] = 10'b1110001000;
mem2[11950] = 10'b1110001000;
mem2[11951] = 10'b1110001000;
mem2[11952] = 10'b1110001000;
mem2[11953] = 10'b1110001000;
mem2[11954] = 10'b1110001000;
mem2[11955] = 10'b1110001000;
mem2[11956] = 10'b1110001000;
mem2[11957] = 10'b1110001000;
mem2[11958] = 10'b1110001001;
mem2[11959] = 10'b1110001001;
mem2[11960] = 10'b1110001001;
mem2[11961] = 10'b1110001001;
mem2[11962] = 10'b1110001001;
mem2[11963] = 10'b1110001001;
mem2[11964] = 10'b1110001001;
mem2[11965] = 10'b1110001001;
mem2[11966] = 10'b1110001001;
mem2[11967] = 10'b1110001001;
mem2[11968] = 10'b1110001001;
mem2[11969] = 10'b1110001001;
mem2[11970] = 10'b1110001001;
mem2[11971] = 10'b1110001001;
mem2[11972] = 10'b1110001001;
mem2[11973] = 10'b1110001010;
mem2[11974] = 10'b1110001010;
mem2[11975] = 10'b1110001010;
mem2[11976] = 10'b1110001010;
mem2[11977] = 10'b1110001010;
mem2[11978] = 10'b1110001010;
mem2[11979] = 10'b1110001010;
mem2[11980] = 10'b1110001010;
mem2[11981] = 10'b1110001010;
mem2[11982] = 10'b1110001010;
mem2[11983] = 10'b1110001010;
mem2[11984] = 10'b1110001010;
mem2[11985] = 10'b1110001010;
mem2[11986] = 10'b1110001010;
mem2[11987] = 10'b1110001010;
mem2[11988] = 10'b1110001011;
mem2[11989] = 10'b1110001011;
mem2[11990] = 10'b1110001011;
mem2[11991] = 10'b1110001011;
mem2[11992] = 10'b1110001011;
mem2[11993] = 10'b1110001011;
mem2[11994] = 10'b1110001011;
mem2[11995] = 10'b1110001011;
mem2[11996] = 10'b1110001011;
mem2[11997] = 10'b1110001011;
mem2[11998] = 10'b1110001011;
mem2[11999] = 10'b1110001011;
mem2[12000] = 10'b1110001011;
mem2[12001] = 10'b1110001011;
mem2[12002] = 10'b1110001011;
mem2[12003] = 10'b1110001100;
mem2[12004] = 10'b1110001100;
mem2[12005] = 10'b1110001100;
mem2[12006] = 10'b1110001100;
mem2[12007] = 10'b1110001100;
mem2[12008] = 10'b1110001100;
mem2[12009] = 10'b1110001100;
mem2[12010] = 10'b1110001100;
mem2[12011] = 10'b1110001100;
mem2[12012] = 10'b1110001100;
mem2[12013] = 10'b1110001100;
mem2[12014] = 10'b1110001100;
mem2[12015] = 10'b1110001100;
mem2[12016] = 10'b1110001100;
mem2[12017] = 10'b1110001100;
mem2[12018] = 10'b1110001101;
mem2[12019] = 10'b1110001101;
mem2[12020] = 10'b1110001101;
mem2[12021] = 10'b1110001101;
mem2[12022] = 10'b1110001101;
mem2[12023] = 10'b1110001101;
mem2[12024] = 10'b1110001101;
mem2[12025] = 10'b1110001101;
mem2[12026] = 10'b1110001101;
mem2[12027] = 10'b1110001101;
mem2[12028] = 10'b1110001101;
mem2[12029] = 10'b1110001101;
mem2[12030] = 10'b1110001101;
mem2[12031] = 10'b1110001101;
mem2[12032] = 10'b1110001101;
mem2[12033] = 10'b1110001110;
mem2[12034] = 10'b1110001110;
mem2[12035] = 10'b1110001110;
mem2[12036] = 10'b1110001110;
mem2[12037] = 10'b1110001110;
mem2[12038] = 10'b1110001110;
mem2[12039] = 10'b1110001110;
mem2[12040] = 10'b1110001110;
mem2[12041] = 10'b1110001110;
mem2[12042] = 10'b1110001110;
mem2[12043] = 10'b1110001110;
mem2[12044] = 10'b1110001110;
mem2[12045] = 10'b1110001110;
mem2[12046] = 10'b1110001110;
mem2[12047] = 10'b1110001110;
mem2[12048] = 10'b1110001110;
mem2[12049] = 10'b1110001111;
mem2[12050] = 10'b1110001111;
mem2[12051] = 10'b1110001111;
mem2[12052] = 10'b1110001111;
mem2[12053] = 10'b1110001111;
mem2[12054] = 10'b1110001111;
mem2[12055] = 10'b1110001111;
mem2[12056] = 10'b1110001111;
mem2[12057] = 10'b1110001111;
mem2[12058] = 10'b1110001111;
mem2[12059] = 10'b1110001111;
mem2[12060] = 10'b1110001111;
mem2[12061] = 10'b1110001111;
mem2[12062] = 10'b1110001111;
mem2[12063] = 10'b1110001111;
mem2[12064] = 10'b1110010000;
mem2[12065] = 10'b1110010000;
mem2[12066] = 10'b1110010000;
mem2[12067] = 10'b1110010000;
mem2[12068] = 10'b1110010000;
mem2[12069] = 10'b1110010000;
mem2[12070] = 10'b1110010000;
mem2[12071] = 10'b1110010000;
mem2[12072] = 10'b1110010000;
mem2[12073] = 10'b1110010000;
mem2[12074] = 10'b1110010000;
mem2[12075] = 10'b1110010000;
mem2[12076] = 10'b1110010000;
mem2[12077] = 10'b1110010000;
mem2[12078] = 10'b1110010000;
mem2[12079] = 10'b1110010001;
mem2[12080] = 10'b1110010001;
mem2[12081] = 10'b1110010001;
mem2[12082] = 10'b1110010001;
mem2[12083] = 10'b1110010001;
mem2[12084] = 10'b1110010001;
mem2[12085] = 10'b1110010001;
mem2[12086] = 10'b1110010001;
mem2[12087] = 10'b1110010001;
mem2[12088] = 10'b1110010001;
mem2[12089] = 10'b1110010001;
mem2[12090] = 10'b1110010001;
mem2[12091] = 10'b1110010001;
mem2[12092] = 10'b1110010001;
mem2[12093] = 10'b1110010001;
mem2[12094] = 10'b1110010001;
mem2[12095] = 10'b1110010010;
mem2[12096] = 10'b1110010010;
mem2[12097] = 10'b1110010010;
mem2[12098] = 10'b1110010010;
mem2[12099] = 10'b1110010010;
mem2[12100] = 10'b1110010010;
mem2[12101] = 10'b1110010010;
mem2[12102] = 10'b1110010010;
mem2[12103] = 10'b1110010010;
mem2[12104] = 10'b1110010010;
mem2[12105] = 10'b1110010010;
mem2[12106] = 10'b1110010010;
mem2[12107] = 10'b1110010010;
mem2[12108] = 10'b1110010010;
mem2[12109] = 10'b1110010010;
mem2[12110] = 10'b1110010011;
mem2[12111] = 10'b1110010011;
mem2[12112] = 10'b1110010011;
mem2[12113] = 10'b1110010011;
mem2[12114] = 10'b1110010011;
mem2[12115] = 10'b1110010011;
mem2[12116] = 10'b1110010011;
mem2[12117] = 10'b1110010011;
mem2[12118] = 10'b1110010011;
mem2[12119] = 10'b1110010011;
mem2[12120] = 10'b1110010011;
mem2[12121] = 10'b1110010011;
mem2[12122] = 10'b1110010011;
mem2[12123] = 10'b1110010011;
mem2[12124] = 10'b1110010011;
mem2[12125] = 10'b1110010011;
mem2[12126] = 10'b1110010100;
mem2[12127] = 10'b1110010100;
mem2[12128] = 10'b1110010100;
mem2[12129] = 10'b1110010100;
mem2[12130] = 10'b1110010100;
mem2[12131] = 10'b1110010100;
mem2[12132] = 10'b1110010100;
mem2[12133] = 10'b1110010100;
mem2[12134] = 10'b1110010100;
mem2[12135] = 10'b1110010100;
mem2[12136] = 10'b1110010100;
mem2[12137] = 10'b1110010100;
mem2[12138] = 10'b1110010100;
mem2[12139] = 10'b1110010100;
mem2[12140] = 10'b1110010100;
mem2[12141] = 10'b1110010101;
mem2[12142] = 10'b1110010101;
mem2[12143] = 10'b1110010101;
mem2[12144] = 10'b1110010101;
mem2[12145] = 10'b1110010101;
mem2[12146] = 10'b1110010101;
mem2[12147] = 10'b1110010101;
mem2[12148] = 10'b1110010101;
mem2[12149] = 10'b1110010101;
mem2[12150] = 10'b1110010101;
mem2[12151] = 10'b1110010101;
mem2[12152] = 10'b1110010101;
mem2[12153] = 10'b1110010101;
mem2[12154] = 10'b1110010101;
mem2[12155] = 10'b1110010101;
mem2[12156] = 10'b1110010101;
mem2[12157] = 10'b1110010110;
mem2[12158] = 10'b1110010110;
mem2[12159] = 10'b1110010110;
mem2[12160] = 10'b1110010110;
mem2[12161] = 10'b1110010110;
mem2[12162] = 10'b1110010110;
mem2[12163] = 10'b1110010110;
mem2[12164] = 10'b1110010110;
mem2[12165] = 10'b1110010110;
mem2[12166] = 10'b1110010110;
mem2[12167] = 10'b1110010110;
mem2[12168] = 10'b1110010110;
mem2[12169] = 10'b1110010110;
mem2[12170] = 10'b1110010110;
mem2[12171] = 10'b1110010110;
mem2[12172] = 10'b1110010111;
mem2[12173] = 10'b1110010111;
mem2[12174] = 10'b1110010111;
mem2[12175] = 10'b1110010111;
mem2[12176] = 10'b1110010111;
mem2[12177] = 10'b1110010111;
mem2[12178] = 10'b1110010111;
mem2[12179] = 10'b1110010111;
mem2[12180] = 10'b1110010111;
mem2[12181] = 10'b1110010111;
mem2[12182] = 10'b1110010111;
mem2[12183] = 10'b1110010111;
mem2[12184] = 10'b1110010111;
mem2[12185] = 10'b1110010111;
mem2[12186] = 10'b1110010111;
mem2[12187] = 10'b1110010111;
mem2[12188] = 10'b1110011000;
mem2[12189] = 10'b1110011000;
mem2[12190] = 10'b1110011000;
mem2[12191] = 10'b1110011000;
mem2[12192] = 10'b1110011000;
mem2[12193] = 10'b1110011000;
mem2[12194] = 10'b1110011000;
mem2[12195] = 10'b1110011000;
mem2[12196] = 10'b1110011000;
mem2[12197] = 10'b1110011000;
mem2[12198] = 10'b1110011000;
mem2[12199] = 10'b1110011000;
mem2[12200] = 10'b1110011000;
mem2[12201] = 10'b1110011000;
mem2[12202] = 10'b1110011000;
mem2[12203] = 10'b1110011000;
mem2[12204] = 10'b1110011001;
mem2[12205] = 10'b1110011001;
mem2[12206] = 10'b1110011001;
mem2[12207] = 10'b1110011001;
mem2[12208] = 10'b1110011001;
mem2[12209] = 10'b1110011001;
mem2[12210] = 10'b1110011001;
mem2[12211] = 10'b1110011001;
mem2[12212] = 10'b1110011001;
mem2[12213] = 10'b1110011001;
mem2[12214] = 10'b1110011001;
mem2[12215] = 10'b1110011001;
mem2[12216] = 10'b1110011001;
mem2[12217] = 10'b1110011001;
mem2[12218] = 10'b1110011001;
mem2[12219] = 10'b1110011001;
mem2[12220] = 10'b1110011010;
mem2[12221] = 10'b1110011010;
mem2[12222] = 10'b1110011010;
mem2[12223] = 10'b1110011010;
mem2[12224] = 10'b1110011010;
mem2[12225] = 10'b1110011010;
mem2[12226] = 10'b1110011010;
mem2[12227] = 10'b1110011010;
mem2[12228] = 10'b1110011010;
mem2[12229] = 10'b1110011010;
mem2[12230] = 10'b1110011010;
mem2[12231] = 10'b1110011010;
mem2[12232] = 10'b1110011010;
mem2[12233] = 10'b1110011010;
mem2[12234] = 10'b1110011010;
mem2[12235] = 10'b1110011010;
mem2[12236] = 10'b1110011011;
mem2[12237] = 10'b1110011011;
mem2[12238] = 10'b1110011011;
mem2[12239] = 10'b1110011011;
mem2[12240] = 10'b1110011011;
mem2[12241] = 10'b1110011011;
mem2[12242] = 10'b1110011011;
mem2[12243] = 10'b1110011011;
mem2[12244] = 10'b1110011011;
mem2[12245] = 10'b1110011011;
mem2[12246] = 10'b1110011011;
mem2[12247] = 10'b1110011011;
mem2[12248] = 10'b1110011011;
mem2[12249] = 10'b1110011011;
mem2[12250] = 10'b1110011011;
mem2[12251] = 10'b1110011011;
mem2[12252] = 10'b1110011100;
mem2[12253] = 10'b1110011100;
mem2[12254] = 10'b1110011100;
mem2[12255] = 10'b1110011100;
mem2[12256] = 10'b1110011100;
mem2[12257] = 10'b1110011100;
mem2[12258] = 10'b1110011100;
mem2[12259] = 10'b1110011100;
mem2[12260] = 10'b1110011100;
mem2[12261] = 10'b1110011100;
mem2[12262] = 10'b1110011100;
mem2[12263] = 10'b1110011100;
mem2[12264] = 10'b1110011100;
mem2[12265] = 10'b1110011100;
mem2[12266] = 10'b1110011100;
mem2[12267] = 10'b1110011100;
mem2[12268] = 10'b1110011101;
mem2[12269] = 10'b1110011101;
mem2[12270] = 10'b1110011101;
mem2[12271] = 10'b1110011101;
mem2[12272] = 10'b1110011101;
mem2[12273] = 10'b1110011101;
mem2[12274] = 10'b1110011101;
mem2[12275] = 10'b1110011101;
mem2[12276] = 10'b1110011101;
mem2[12277] = 10'b1110011101;
mem2[12278] = 10'b1110011101;
mem2[12279] = 10'b1110011101;
mem2[12280] = 10'b1110011101;
mem2[12281] = 10'b1110011101;
mem2[12282] = 10'b1110011101;
mem2[12283] = 10'b1110011101;
mem2[12284] = 10'b1110011110;
mem2[12285] = 10'b1110011110;
mem2[12286] = 10'b1110011110;
mem2[12287] = 10'b1110011110;
mem2[12288] = 10'b1110011110;
mem2[12289] = 10'b1110011110;
mem2[12290] = 10'b1110011110;
mem2[12291] = 10'b1110011110;
mem2[12292] = 10'b1110011110;
mem2[12293] = 10'b1110011110;
mem2[12294] = 10'b1110011110;
mem2[12295] = 10'b1110011110;
mem2[12296] = 10'b1110011110;
mem2[12297] = 10'b1110011110;
mem2[12298] = 10'b1110011110;
mem2[12299] = 10'b1110011110;
mem2[12300] = 10'b1110011110;
mem2[12301] = 10'b1110011111;
mem2[12302] = 10'b1110011111;
mem2[12303] = 10'b1110011111;
mem2[12304] = 10'b1110011111;
mem2[12305] = 10'b1110011111;
mem2[12306] = 10'b1110011111;
mem2[12307] = 10'b1110011111;
mem2[12308] = 10'b1110011111;
mem2[12309] = 10'b1110011111;
mem2[12310] = 10'b1110011111;
mem2[12311] = 10'b1110011111;
mem2[12312] = 10'b1110011111;
mem2[12313] = 10'b1110011111;
mem2[12314] = 10'b1110011111;
mem2[12315] = 10'b1110011111;
mem2[12316] = 10'b1110011111;
mem2[12317] = 10'b1110100000;
mem2[12318] = 10'b1110100000;
mem2[12319] = 10'b1110100000;
mem2[12320] = 10'b1110100000;
mem2[12321] = 10'b1110100000;
mem2[12322] = 10'b1110100000;
mem2[12323] = 10'b1110100000;
mem2[12324] = 10'b1110100000;
mem2[12325] = 10'b1110100000;
mem2[12326] = 10'b1110100000;
mem2[12327] = 10'b1110100000;
mem2[12328] = 10'b1110100000;
mem2[12329] = 10'b1110100000;
mem2[12330] = 10'b1110100000;
mem2[12331] = 10'b1110100000;
mem2[12332] = 10'b1110100000;
mem2[12333] = 10'b1110100001;
mem2[12334] = 10'b1110100001;
mem2[12335] = 10'b1110100001;
mem2[12336] = 10'b1110100001;
mem2[12337] = 10'b1110100001;
mem2[12338] = 10'b1110100001;
mem2[12339] = 10'b1110100001;
mem2[12340] = 10'b1110100001;
mem2[12341] = 10'b1110100001;
mem2[12342] = 10'b1110100001;
mem2[12343] = 10'b1110100001;
mem2[12344] = 10'b1110100001;
mem2[12345] = 10'b1110100001;
mem2[12346] = 10'b1110100001;
mem2[12347] = 10'b1110100001;
mem2[12348] = 10'b1110100001;
mem2[12349] = 10'b1110100001;
mem2[12350] = 10'b1110100010;
mem2[12351] = 10'b1110100010;
mem2[12352] = 10'b1110100010;
mem2[12353] = 10'b1110100010;
mem2[12354] = 10'b1110100010;
mem2[12355] = 10'b1110100010;
mem2[12356] = 10'b1110100010;
mem2[12357] = 10'b1110100010;
mem2[12358] = 10'b1110100010;
mem2[12359] = 10'b1110100010;
mem2[12360] = 10'b1110100010;
mem2[12361] = 10'b1110100010;
mem2[12362] = 10'b1110100010;
mem2[12363] = 10'b1110100010;
mem2[12364] = 10'b1110100010;
mem2[12365] = 10'b1110100010;
mem2[12366] = 10'b1110100011;
mem2[12367] = 10'b1110100011;
mem2[12368] = 10'b1110100011;
mem2[12369] = 10'b1110100011;
mem2[12370] = 10'b1110100011;
mem2[12371] = 10'b1110100011;
mem2[12372] = 10'b1110100011;
mem2[12373] = 10'b1110100011;
mem2[12374] = 10'b1110100011;
mem2[12375] = 10'b1110100011;
mem2[12376] = 10'b1110100011;
mem2[12377] = 10'b1110100011;
mem2[12378] = 10'b1110100011;
mem2[12379] = 10'b1110100011;
mem2[12380] = 10'b1110100011;
mem2[12381] = 10'b1110100011;
mem2[12382] = 10'b1110100011;
mem2[12383] = 10'b1110100100;
mem2[12384] = 10'b1110100100;
mem2[12385] = 10'b1110100100;
mem2[12386] = 10'b1110100100;
mem2[12387] = 10'b1110100100;
mem2[12388] = 10'b1110100100;
mem2[12389] = 10'b1110100100;
mem2[12390] = 10'b1110100100;
mem2[12391] = 10'b1110100100;
mem2[12392] = 10'b1110100100;
mem2[12393] = 10'b1110100100;
mem2[12394] = 10'b1110100100;
mem2[12395] = 10'b1110100100;
mem2[12396] = 10'b1110100100;
mem2[12397] = 10'b1110100100;
mem2[12398] = 10'b1110100100;
mem2[12399] = 10'b1110100100;
mem2[12400] = 10'b1110100101;
mem2[12401] = 10'b1110100101;
mem2[12402] = 10'b1110100101;
mem2[12403] = 10'b1110100101;
mem2[12404] = 10'b1110100101;
mem2[12405] = 10'b1110100101;
mem2[12406] = 10'b1110100101;
mem2[12407] = 10'b1110100101;
mem2[12408] = 10'b1110100101;
mem2[12409] = 10'b1110100101;
mem2[12410] = 10'b1110100101;
mem2[12411] = 10'b1110100101;
mem2[12412] = 10'b1110100101;
mem2[12413] = 10'b1110100101;
mem2[12414] = 10'b1110100101;
mem2[12415] = 10'b1110100101;
mem2[12416] = 10'b1110100101;
mem2[12417] = 10'b1110100110;
mem2[12418] = 10'b1110100110;
mem2[12419] = 10'b1110100110;
mem2[12420] = 10'b1110100110;
mem2[12421] = 10'b1110100110;
mem2[12422] = 10'b1110100110;
mem2[12423] = 10'b1110100110;
mem2[12424] = 10'b1110100110;
mem2[12425] = 10'b1110100110;
mem2[12426] = 10'b1110100110;
mem2[12427] = 10'b1110100110;
mem2[12428] = 10'b1110100110;
mem2[12429] = 10'b1110100110;
mem2[12430] = 10'b1110100110;
mem2[12431] = 10'b1110100110;
mem2[12432] = 10'b1110100110;
mem2[12433] = 10'b1110100110;
mem2[12434] = 10'b1110100111;
mem2[12435] = 10'b1110100111;
mem2[12436] = 10'b1110100111;
mem2[12437] = 10'b1110100111;
mem2[12438] = 10'b1110100111;
mem2[12439] = 10'b1110100111;
mem2[12440] = 10'b1110100111;
mem2[12441] = 10'b1110100111;
mem2[12442] = 10'b1110100111;
mem2[12443] = 10'b1110100111;
mem2[12444] = 10'b1110100111;
mem2[12445] = 10'b1110100111;
mem2[12446] = 10'b1110100111;
mem2[12447] = 10'b1110100111;
mem2[12448] = 10'b1110100111;
mem2[12449] = 10'b1110100111;
mem2[12450] = 10'b1110100111;
mem2[12451] = 10'b1110101000;
mem2[12452] = 10'b1110101000;
mem2[12453] = 10'b1110101000;
mem2[12454] = 10'b1110101000;
mem2[12455] = 10'b1110101000;
mem2[12456] = 10'b1110101000;
mem2[12457] = 10'b1110101000;
mem2[12458] = 10'b1110101000;
mem2[12459] = 10'b1110101000;
mem2[12460] = 10'b1110101000;
mem2[12461] = 10'b1110101000;
mem2[12462] = 10'b1110101000;
mem2[12463] = 10'b1110101000;
mem2[12464] = 10'b1110101000;
mem2[12465] = 10'b1110101000;
mem2[12466] = 10'b1110101000;
mem2[12467] = 10'b1110101000;
mem2[12468] = 10'b1110101001;
mem2[12469] = 10'b1110101001;
mem2[12470] = 10'b1110101001;
mem2[12471] = 10'b1110101001;
mem2[12472] = 10'b1110101001;
mem2[12473] = 10'b1110101001;
mem2[12474] = 10'b1110101001;
mem2[12475] = 10'b1110101001;
mem2[12476] = 10'b1110101001;
mem2[12477] = 10'b1110101001;
mem2[12478] = 10'b1110101001;
mem2[12479] = 10'b1110101001;
mem2[12480] = 10'b1110101001;
mem2[12481] = 10'b1110101001;
mem2[12482] = 10'b1110101001;
mem2[12483] = 10'b1110101001;
mem2[12484] = 10'b1110101001;
mem2[12485] = 10'b1110101010;
mem2[12486] = 10'b1110101010;
mem2[12487] = 10'b1110101010;
mem2[12488] = 10'b1110101010;
mem2[12489] = 10'b1110101010;
mem2[12490] = 10'b1110101010;
mem2[12491] = 10'b1110101010;
mem2[12492] = 10'b1110101010;
mem2[12493] = 10'b1110101010;
mem2[12494] = 10'b1110101010;
mem2[12495] = 10'b1110101010;
mem2[12496] = 10'b1110101010;
mem2[12497] = 10'b1110101010;
mem2[12498] = 10'b1110101010;
mem2[12499] = 10'b1110101010;
mem2[12500] = 10'b1110101010;
mem2[12501] = 10'b1110101010;
mem2[12502] = 10'b1110101011;
mem2[12503] = 10'b1110101011;
mem2[12504] = 10'b1110101011;
mem2[12505] = 10'b1110101011;
mem2[12506] = 10'b1110101011;
mem2[12507] = 10'b1110101011;
mem2[12508] = 10'b1110101011;
mem2[12509] = 10'b1110101011;
mem2[12510] = 10'b1110101011;
mem2[12511] = 10'b1110101011;
mem2[12512] = 10'b1110101011;
mem2[12513] = 10'b1110101011;
mem2[12514] = 10'b1110101011;
mem2[12515] = 10'b1110101011;
mem2[12516] = 10'b1110101011;
mem2[12517] = 10'b1110101011;
mem2[12518] = 10'b1110101011;
mem2[12519] = 10'b1110101100;
mem2[12520] = 10'b1110101100;
mem2[12521] = 10'b1110101100;
mem2[12522] = 10'b1110101100;
mem2[12523] = 10'b1110101100;
mem2[12524] = 10'b1110101100;
mem2[12525] = 10'b1110101100;
mem2[12526] = 10'b1110101100;
mem2[12527] = 10'b1110101100;
mem2[12528] = 10'b1110101100;
mem2[12529] = 10'b1110101100;
mem2[12530] = 10'b1110101100;
mem2[12531] = 10'b1110101100;
mem2[12532] = 10'b1110101100;
mem2[12533] = 10'b1110101100;
mem2[12534] = 10'b1110101100;
mem2[12535] = 10'b1110101100;
mem2[12536] = 10'b1110101100;
mem2[12537] = 10'b1110101101;
mem2[12538] = 10'b1110101101;
mem2[12539] = 10'b1110101101;
mem2[12540] = 10'b1110101101;
mem2[12541] = 10'b1110101101;
mem2[12542] = 10'b1110101101;
mem2[12543] = 10'b1110101101;
mem2[12544] = 10'b1110101101;
mem2[12545] = 10'b1110101101;
mem2[12546] = 10'b1110101101;
mem2[12547] = 10'b1110101101;
mem2[12548] = 10'b1110101101;
mem2[12549] = 10'b1110101101;
mem2[12550] = 10'b1110101101;
mem2[12551] = 10'b1110101101;
mem2[12552] = 10'b1110101101;
mem2[12553] = 10'b1110101101;
mem2[12554] = 10'b1110101110;
mem2[12555] = 10'b1110101110;
mem2[12556] = 10'b1110101110;
mem2[12557] = 10'b1110101110;
mem2[12558] = 10'b1110101110;
mem2[12559] = 10'b1110101110;
mem2[12560] = 10'b1110101110;
mem2[12561] = 10'b1110101110;
mem2[12562] = 10'b1110101110;
mem2[12563] = 10'b1110101110;
mem2[12564] = 10'b1110101110;
mem2[12565] = 10'b1110101110;
mem2[12566] = 10'b1110101110;
mem2[12567] = 10'b1110101110;
mem2[12568] = 10'b1110101110;
mem2[12569] = 10'b1110101110;
mem2[12570] = 10'b1110101110;
mem2[12571] = 10'b1110101110;
mem2[12572] = 10'b1110101111;
mem2[12573] = 10'b1110101111;
mem2[12574] = 10'b1110101111;
mem2[12575] = 10'b1110101111;
mem2[12576] = 10'b1110101111;
mem2[12577] = 10'b1110101111;
mem2[12578] = 10'b1110101111;
mem2[12579] = 10'b1110101111;
mem2[12580] = 10'b1110101111;
mem2[12581] = 10'b1110101111;
mem2[12582] = 10'b1110101111;
mem2[12583] = 10'b1110101111;
mem2[12584] = 10'b1110101111;
mem2[12585] = 10'b1110101111;
mem2[12586] = 10'b1110101111;
mem2[12587] = 10'b1110101111;
mem2[12588] = 10'b1110101111;
mem2[12589] = 10'b1110101111;
mem2[12590] = 10'b1110110000;
mem2[12591] = 10'b1110110000;
mem2[12592] = 10'b1110110000;
mem2[12593] = 10'b1110110000;
mem2[12594] = 10'b1110110000;
mem2[12595] = 10'b1110110000;
mem2[12596] = 10'b1110110000;
mem2[12597] = 10'b1110110000;
mem2[12598] = 10'b1110110000;
mem2[12599] = 10'b1110110000;
mem2[12600] = 10'b1110110000;
mem2[12601] = 10'b1110110000;
mem2[12602] = 10'b1110110000;
mem2[12603] = 10'b1110110000;
mem2[12604] = 10'b1110110000;
mem2[12605] = 10'b1110110000;
mem2[12606] = 10'b1110110000;
mem2[12607] = 10'b1110110000;
mem2[12608] = 10'b1110110001;
mem2[12609] = 10'b1110110001;
mem2[12610] = 10'b1110110001;
mem2[12611] = 10'b1110110001;
mem2[12612] = 10'b1110110001;
mem2[12613] = 10'b1110110001;
mem2[12614] = 10'b1110110001;
mem2[12615] = 10'b1110110001;
mem2[12616] = 10'b1110110001;
mem2[12617] = 10'b1110110001;
mem2[12618] = 10'b1110110001;
mem2[12619] = 10'b1110110001;
mem2[12620] = 10'b1110110001;
mem2[12621] = 10'b1110110001;
mem2[12622] = 10'b1110110001;
mem2[12623] = 10'b1110110001;
mem2[12624] = 10'b1110110001;
mem2[12625] = 10'b1110110001;
mem2[12626] = 10'b1110110010;
mem2[12627] = 10'b1110110010;
mem2[12628] = 10'b1110110010;
mem2[12629] = 10'b1110110010;
mem2[12630] = 10'b1110110010;
mem2[12631] = 10'b1110110010;
mem2[12632] = 10'b1110110010;
mem2[12633] = 10'b1110110010;
mem2[12634] = 10'b1110110010;
mem2[12635] = 10'b1110110010;
mem2[12636] = 10'b1110110010;
mem2[12637] = 10'b1110110010;
mem2[12638] = 10'b1110110010;
mem2[12639] = 10'b1110110010;
mem2[12640] = 10'b1110110010;
mem2[12641] = 10'b1110110010;
mem2[12642] = 10'b1110110010;
mem2[12643] = 10'b1110110010;
mem2[12644] = 10'b1110110011;
mem2[12645] = 10'b1110110011;
mem2[12646] = 10'b1110110011;
mem2[12647] = 10'b1110110011;
mem2[12648] = 10'b1110110011;
mem2[12649] = 10'b1110110011;
mem2[12650] = 10'b1110110011;
mem2[12651] = 10'b1110110011;
mem2[12652] = 10'b1110110011;
mem2[12653] = 10'b1110110011;
mem2[12654] = 10'b1110110011;
mem2[12655] = 10'b1110110011;
mem2[12656] = 10'b1110110011;
mem2[12657] = 10'b1110110011;
mem2[12658] = 10'b1110110011;
mem2[12659] = 10'b1110110011;
mem2[12660] = 10'b1110110011;
mem2[12661] = 10'b1110110011;
mem2[12662] = 10'b1110110100;
mem2[12663] = 10'b1110110100;
mem2[12664] = 10'b1110110100;
mem2[12665] = 10'b1110110100;
mem2[12666] = 10'b1110110100;
mem2[12667] = 10'b1110110100;
mem2[12668] = 10'b1110110100;
mem2[12669] = 10'b1110110100;
mem2[12670] = 10'b1110110100;
mem2[12671] = 10'b1110110100;
mem2[12672] = 10'b1110110100;
mem2[12673] = 10'b1110110100;
mem2[12674] = 10'b1110110100;
mem2[12675] = 10'b1110110100;
mem2[12676] = 10'b1110110100;
mem2[12677] = 10'b1110110100;
mem2[12678] = 10'b1110110100;
mem2[12679] = 10'b1110110100;
mem2[12680] = 10'b1110110101;
mem2[12681] = 10'b1110110101;
mem2[12682] = 10'b1110110101;
mem2[12683] = 10'b1110110101;
mem2[12684] = 10'b1110110101;
mem2[12685] = 10'b1110110101;
mem2[12686] = 10'b1110110101;
mem2[12687] = 10'b1110110101;
mem2[12688] = 10'b1110110101;
mem2[12689] = 10'b1110110101;
mem2[12690] = 10'b1110110101;
mem2[12691] = 10'b1110110101;
mem2[12692] = 10'b1110110101;
mem2[12693] = 10'b1110110101;
mem2[12694] = 10'b1110110101;
mem2[12695] = 10'b1110110101;
mem2[12696] = 10'b1110110101;
mem2[12697] = 10'b1110110101;
mem2[12698] = 10'b1110110110;
mem2[12699] = 10'b1110110110;
mem2[12700] = 10'b1110110110;
mem2[12701] = 10'b1110110110;
mem2[12702] = 10'b1110110110;
mem2[12703] = 10'b1110110110;
mem2[12704] = 10'b1110110110;
mem2[12705] = 10'b1110110110;
mem2[12706] = 10'b1110110110;
mem2[12707] = 10'b1110110110;
mem2[12708] = 10'b1110110110;
mem2[12709] = 10'b1110110110;
mem2[12710] = 10'b1110110110;
mem2[12711] = 10'b1110110110;
mem2[12712] = 10'b1110110110;
mem2[12713] = 10'b1110110110;
mem2[12714] = 10'b1110110110;
mem2[12715] = 10'b1110110110;
mem2[12716] = 10'b1110110110;
mem2[12717] = 10'b1110110111;
mem2[12718] = 10'b1110110111;
mem2[12719] = 10'b1110110111;
mem2[12720] = 10'b1110110111;
mem2[12721] = 10'b1110110111;
mem2[12722] = 10'b1110110111;
mem2[12723] = 10'b1110110111;
mem2[12724] = 10'b1110110111;
mem2[12725] = 10'b1110110111;
mem2[12726] = 10'b1110110111;
mem2[12727] = 10'b1110110111;
mem2[12728] = 10'b1110110111;
mem2[12729] = 10'b1110110111;
mem2[12730] = 10'b1110110111;
mem2[12731] = 10'b1110110111;
mem2[12732] = 10'b1110110111;
mem2[12733] = 10'b1110110111;
mem2[12734] = 10'b1110110111;
mem2[12735] = 10'b1110110111;
mem2[12736] = 10'b1110111000;
mem2[12737] = 10'b1110111000;
mem2[12738] = 10'b1110111000;
mem2[12739] = 10'b1110111000;
mem2[12740] = 10'b1110111000;
mem2[12741] = 10'b1110111000;
mem2[12742] = 10'b1110111000;
mem2[12743] = 10'b1110111000;
mem2[12744] = 10'b1110111000;
mem2[12745] = 10'b1110111000;
mem2[12746] = 10'b1110111000;
mem2[12747] = 10'b1110111000;
mem2[12748] = 10'b1110111000;
mem2[12749] = 10'b1110111000;
mem2[12750] = 10'b1110111000;
mem2[12751] = 10'b1110111000;
mem2[12752] = 10'b1110111000;
mem2[12753] = 10'b1110111000;
mem2[12754] = 10'b1110111001;
mem2[12755] = 10'b1110111001;
mem2[12756] = 10'b1110111001;
mem2[12757] = 10'b1110111001;
mem2[12758] = 10'b1110111001;
mem2[12759] = 10'b1110111001;
mem2[12760] = 10'b1110111001;
mem2[12761] = 10'b1110111001;
mem2[12762] = 10'b1110111001;
mem2[12763] = 10'b1110111001;
mem2[12764] = 10'b1110111001;
mem2[12765] = 10'b1110111001;
mem2[12766] = 10'b1110111001;
mem2[12767] = 10'b1110111001;
mem2[12768] = 10'b1110111001;
mem2[12769] = 10'b1110111001;
mem2[12770] = 10'b1110111001;
mem2[12771] = 10'b1110111001;
mem2[12772] = 10'b1110111001;
mem2[12773] = 10'b1110111010;
mem2[12774] = 10'b1110111010;
mem2[12775] = 10'b1110111010;
mem2[12776] = 10'b1110111010;
mem2[12777] = 10'b1110111010;
mem2[12778] = 10'b1110111010;
mem2[12779] = 10'b1110111010;
mem2[12780] = 10'b1110111010;
mem2[12781] = 10'b1110111010;
mem2[12782] = 10'b1110111010;
mem2[12783] = 10'b1110111010;
mem2[12784] = 10'b1110111010;
mem2[12785] = 10'b1110111010;
mem2[12786] = 10'b1110111010;
mem2[12787] = 10'b1110111010;
mem2[12788] = 10'b1110111010;
mem2[12789] = 10'b1110111010;
mem2[12790] = 10'b1110111010;
mem2[12791] = 10'b1110111010;
mem2[12792] = 10'b1110111011;
mem2[12793] = 10'b1110111011;
mem2[12794] = 10'b1110111011;
mem2[12795] = 10'b1110111011;
mem2[12796] = 10'b1110111011;
mem2[12797] = 10'b1110111011;
mem2[12798] = 10'b1110111011;
mem2[12799] = 10'b1110111011;
mem2[12800] = 10'b1110111011;
mem2[12801] = 10'b1110111011;
mem2[12802] = 10'b1110111011;
mem2[12803] = 10'b1110111011;
mem2[12804] = 10'b1110111011;
mem2[12805] = 10'b1110111011;
mem2[12806] = 10'b1110111011;
mem2[12807] = 10'b1110111011;
mem2[12808] = 10'b1110111011;
mem2[12809] = 10'b1110111011;
mem2[12810] = 10'b1110111011;
mem2[12811] = 10'b1110111100;
mem2[12812] = 10'b1110111100;
mem2[12813] = 10'b1110111100;
mem2[12814] = 10'b1110111100;
mem2[12815] = 10'b1110111100;
mem2[12816] = 10'b1110111100;
mem2[12817] = 10'b1110111100;
mem2[12818] = 10'b1110111100;
mem2[12819] = 10'b1110111100;
mem2[12820] = 10'b1110111100;
mem2[12821] = 10'b1110111100;
mem2[12822] = 10'b1110111100;
mem2[12823] = 10'b1110111100;
mem2[12824] = 10'b1110111100;
mem2[12825] = 10'b1110111100;
mem2[12826] = 10'b1110111100;
mem2[12827] = 10'b1110111100;
mem2[12828] = 10'b1110111100;
mem2[12829] = 10'b1110111100;
mem2[12830] = 10'b1110111101;
mem2[12831] = 10'b1110111101;
mem2[12832] = 10'b1110111101;
mem2[12833] = 10'b1110111101;
mem2[12834] = 10'b1110111101;
mem2[12835] = 10'b1110111101;
mem2[12836] = 10'b1110111101;
mem2[12837] = 10'b1110111101;
mem2[12838] = 10'b1110111101;
mem2[12839] = 10'b1110111101;
mem2[12840] = 10'b1110111101;
mem2[12841] = 10'b1110111101;
mem2[12842] = 10'b1110111101;
mem2[12843] = 10'b1110111101;
mem2[12844] = 10'b1110111101;
mem2[12845] = 10'b1110111101;
mem2[12846] = 10'b1110111101;
mem2[12847] = 10'b1110111101;
mem2[12848] = 10'b1110111101;
mem2[12849] = 10'b1110111101;
mem2[12850] = 10'b1110111110;
mem2[12851] = 10'b1110111110;
mem2[12852] = 10'b1110111110;
mem2[12853] = 10'b1110111110;
mem2[12854] = 10'b1110111110;
mem2[12855] = 10'b1110111110;
mem2[12856] = 10'b1110111110;
mem2[12857] = 10'b1110111110;
mem2[12858] = 10'b1110111110;
mem2[12859] = 10'b1110111110;
mem2[12860] = 10'b1110111110;
mem2[12861] = 10'b1110111110;
mem2[12862] = 10'b1110111110;
mem2[12863] = 10'b1110111110;
mem2[12864] = 10'b1110111110;
mem2[12865] = 10'b1110111110;
mem2[12866] = 10'b1110111110;
mem2[12867] = 10'b1110111110;
mem2[12868] = 10'b1110111110;
mem2[12869] = 10'b1110111111;
mem2[12870] = 10'b1110111111;
mem2[12871] = 10'b1110111111;
mem2[12872] = 10'b1110111111;
mem2[12873] = 10'b1110111111;
mem2[12874] = 10'b1110111111;
mem2[12875] = 10'b1110111111;
mem2[12876] = 10'b1110111111;
mem2[12877] = 10'b1110111111;
mem2[12878] = 10'b1110111111;
mem2[12879] = 10'b1110111111;
mem2[12880] = 10'b1110111111;
mem2[12881] = 10'b1110111111;
mem2[12882] = 10'b1110111111;
mem2[12883] = 10'b1110111111;
mem2[12884] = 10'b1110111111;
mem2[12885] = 10'b1110111111;
mem2[12886] = 10'b1110111111;
mem2[12887] = 10'b1110111111;
mem2[12888] = 10'b1110111111;
mem2[12889] = 10'b1111000000;
mem2[12890] = 10'b1111000000;
mem2[12891] = 10'b1111000000;
mem2[12892] = 10'b1111000000;
mem2[12893] = 10'b1111000000;
mem2[12894] = 10'b1111000000;
mem2[12895] = 10'b1111000000;
mem2[12896] = 10'b1111000000;
mem2[12897] = 10'b1111000000;
mem2[12898] = 10'b1111000000;
mem2[12899] = 10'b1111000000;
mem2[12900] = 10'b1111000000;
mem2[12901] = 10'b1111000000;
mem2[12902] = 10'b1111000000;
mem2[12903] = 10'b1111000000;
mem2[12904] = 10'b1111000000;
mem2[12905] = 10'b1111000000;
mem2[12906] = 10'b1111000000;
mem2[12907] = 10'b1111000000;
mem2[12908] = 10'b1111000000;
mem2[12909] = 10'b1111000001;
mem2[12910] = 10'b1111000001;
mem2[12911] = 10'b1111000001;
mem2[12912] = 10'b1111000001;
mem2[12913] = 10'b1111000001;
mem2[12914] = 10'b1111000001;
mem2[12915] = 10'b1111000001;
mem2[12916] = 10'b1111000001;
mem2[12917] = 10'b1111000001;
mem2[12918] = 10'b1111000001;
mem2[12919] = 10'b1111000001;
mem2[12920] = 10'b1111000001;
mem2[12921] = 10'b1111000001;
mem2[12922] = 10'b1111000001;
mem2[12923] = 10'b1111000001;
mem2[12924] = 10'b1111000001;
mem2[12925] = 10'b1111000001;
mem2[12926] = 10'b1111000001;
mem2[12927] = 10'b1111000001;
mem2[12928] = 10'b1111000001;
mem2[12929] = 10'b1111000010;
mem2[12930] = 10'b1111000010;
mem2[12931] = 10'b1111000010;
mem2[12932] = 10'b1111000010;
mem2[12933] = 10'b1111000010;
mem2[12934] = 10'b1111000010;
mem2[12935] = 10'b1111000010;
mem2[12936] = 10'b1111000010;
mem2[12937] = 10'b1111000010;
mem2[12938] = 10'b1111000010;
mem2[12939] = 10'b1111000010;
mem2[12940] = 10'b1111000010;
mem2[12941] = 10'b1111000010;
mem2[12942] = 10'b1111000010;
mem2[12943] = 10'b1111000010;
mem2[12944] = 10'b1111000010;
mem2[12945] = 10'b1111000010;
mem2[12946] = 10'b1111000010;
mem2[12947] = 10'b1111000010;
mem2[12948] = 10'b1111000010;
mem2[12949] = 10'b1111000011;
mem2[12950] = 10'b1111000011;
mem2[12951] = 10'b1111000011;
mem2[12952] = 10'b1111000011;
mem2[12953] = 10'b1111000011;
mem2[12954] = 10'b1111000011;
mem2[12955] = 10'b1111000011;
mem2[12956] = 10'b1111000011;
mem2[12957] = 10'b1111000011;
mem2[12958] = 10'b1111000011;
mem2[12959] = 10'b1111000011;
mem2[12960] = 10'b1111000011;
mem2[12961] = 10'b1111000011;
mem2[12962] = 10'b1111000011;
mem2[12963] = 10'b1111000011;
mem2[12964] = 10'b1111000011;
mem2[12965] = 10'b1111000011;
mem2[12966] = 10'b1111000011;
mem2[12967] = 10'b1111000011;
mem2[12968] = 10'b1111000011;
mem2[12969] = 10'b1111000100;
mem2[12970] = 10'b1111000100;
mem2[12971] = 10'b1111000100;
mem2[12972] = 10'b1111000100;
mem2[12973] = 10'b1111000100;
mem2[12974] = 10'b1111000100;
mem2[12975] = 10'b1111000100;
mem2[12976] = 10'b1111000100;
mem2[12977] = 10'b1111000100;
mem2[12978] = 10'b1111000100;
mem2[12979] = 10'b1111000100;
mem2[12980] = 10'b1111000100;
mem2[12981] = 10'b1111000100;
mem2[12982] = 10'b1111000100;
mem2[12983] = 10'b1111000100;
mem2[12984] = 10'b1111000100;
mem2[12985] = 10'b1111000100;
mem2[12986] = 10'b1111000100;
mem2[12987] = 10'b1111000100;
mem2[12988] = 10'b1111000100;
mem2[12989] = 10'b1111000101;
mem2[12990] = 10'b1111000101;
mem2[12991] = 10'b1111000101;
mem2[12992] = 10'b1111000101;
mem2[12993] = 10'b1111000101;
mem2[12994] = 10'b1111000101;
mem2[12995] = 10'b1111000101;
mem2[12996] = 10'b1111000101;
mem2[12997] = 10'b1111000101;
mem2[12998] = 10'b1111000101;
mem2[12999] = 10'b1111000101;
mem2[13000] = 10'b1111000101;
mem2[13001] = 10'b1111000101;
mem2[13002] = 10'b1111000101;
mem2[13003] = 10'b1111000101;
mem2[13004] = 10'b1111000101;
mem2[13005] = 10'b1111000101;
mem2[13006] = 10'b1111000101;
mem2[13007] = 10'b1111000101;
mem2[13008] = 10'b1111000101;
mem2[13009] = 10'b1111000101;
mem2[13010] = 10'b1111000110;
mem2[13011] = 10'b1111000110;
mem2[13012] = 10'b1111000110;
mem2[13013] = 10'b1111000110;
mem2[13014] = 10'b1111000110;
mem2[13015] = 10'b1111000110;
mem2[13016] = 10'b1111000110;
mem2[13017] = 10'b1111000110;
mem2[13018] = 10'b1111000110;
mem2[13019] = 10'b1111000110;
mem2[13020] = 10'b1111000110;
mem2[13021] = 10'b1111000110;
mem2[13022] = 10'b1111000110;
mem2[13023] = 10'b1111000110;
mem2[13024] = 10'b1111000110;
mem2[13025] = 10'b1111000110;
mem2[13026] = 10'b1111000110;
mem2[13027] = 10'b1111000110;
mem2[13028] = 10'b1111000110;
mem2[13029] = 10'b1111000110;
mem2[13030] = 10'b1111000110;
mem2[13031] = 10'b1111000111;
mem2[13032] = 10'b1111000111;
mem2[13033] = 10'b1111000111;
mem2[13034] = 10'b1111000111;
mem2[13035] = 10'b1111000111;
mem2[13036] = 10'b1111000111;
mem2[13037] = 10'b1111000111;
mem2[13038] = 10'b1111000111;
mem2[13039] = 10'b1111000111;
mem2[13040] = 10'b1111000111;
mem2[13041] = 10'b1111000111;
mem2[13042] = 10'b1111000111;
mem2[13043] = 10'b1111000111;
mem2[13044] = 10'b1111000111;
mem2[13045] = 10'b1111000111;
mem2[13046] = 10'b1111000111;
mem2[13047] = 10'b1111000111;
mem2[13048] = 10'b1111000111;
mem2[13049] = 10'b1111000111;
mem2[13050] = 10'b1111000111;
mem2[13051] = 10'b1111000111;
mem2[13052] = 10'b1111001000;
mem2[13053] = 10'b1111001000;
mem2[13054] = 10'b1111001000;
mem2[13055] = 10'b1111001000;
mem2[13056] = 10'b1111001000;
mem2[13057] = 10'b1111001000;
mem2[13058] = 10'b1111001000;
mem2[13059] = 10'b1111001000;
mem2[13060] = 10'b1111001000;
mem2[13061] = 10'b1111001000;
mem2[13062] = 10'b1111001000;
mem2[13063] = 10'b1111001000;
mem2[13064] = 10'b1111001000;
mem2[13065] = 10'b1111001000;
mem2[13066] = 10'b1111001000;
mem2[13067] = 10'b1111001000;
mem2[13068] = 10'b1111001000;
mem2[13069] = 10'b1111001000;
mem2[13070] = 10'b1111001000;
mem2[13071] = 10'b1111001000;
mem2[13072] = 10'b1111001000;
mem2[13073] = 10'b1111001001;
mem2[13074] = 10'b1111001001;
mem2[13075] = 10'b1111001001;
mem2[13076] = 10'b1111001001;
mem2[13077] = 10'b1111001001;
mem2[13078] = 10'b1111001001;
mem2[13079] = 10'b1111001001;
mem2[13080] = 10'b1111001001;
mem2[13081] = 10'b1111001001;
mem2[13082] = 10'b1111001001;
mem2[13083] = 10'b1111001001;
mem2[13084] = 10'b1111001001;
mem2[13085] = 10'b1111001001;
mem2[13086] = 10'b1111001001;
mem2[13087] = 10'b1111001001;
mem2[13088] = 10'b1111001001;
mem2[13089] = 10'b1111001001;
mem2[13090] = 10'b1111001001;
mem2[13091] = 10'b1111001001;
mem2[13092] = 10'b1111001001;
mem2[13093] = 10'b1111001001;
mem2[13094] = 10'b1111001010;
mem2[13095] = 10'b1111001010;
mem2[13096] = 10'b1111001010;
mem2[13097] = 10'b1111001010;
mem2[13098] = 10'b1111001010;
mem2[13099] = 10'b1111001010;
mem2[13100] = 10'b1111001010;
mem2[13101] = 10'b1111001010;
mem2[13102] = 10'b1111001010;
mem2[13103] = 10'b1111001010;
mem2[13104] = 10'b1111001010;
mem2[13105] = 10'b1111001010;
mem2[13106] = 10'b1111001010;
mem2[13107] = 10'b1111001010;
mem2[13108] = 10'b1111001010;
mem2[13109] = 10'b1111001010;
mem2[13110] = 10'b1111001010;
mem2[13111] = 10'b1111001010;
mem2[13112] = 10'b1111001010;
mem2[13113] = 10'b1111001010;
mem2[13114] = 10'b1111001010;
mem2[13115] = 10'b1111001010;
mem2[13116] = 10'b1111001011;
mem2[13117] = 10'b1111001011;
mem2[13118] = 10'b1111001011;
mem2[13119] = 10'b1111001011;
mem2[13120] = 10'b1111001011;
mem2[13121] = 10'b1111001011;
mem2[13122] = 10'b1111001011;
mem2[13123] = 10'b1111001011;
mem2[13124] = 10'b1111001011;
mem2[13125] = 10'b1111001011;
mem2[13126] = 10'b1111001011;
mem2[13127] = 10'b1111001011;
mem2[13128] = 10'b1111001011;
mem2[13129] = 10'b1111001011;
mem2[13130] = 10'b1111001011;
mem2[13131] = 10'b1111001011;
mem2[13132] = 10'b1111001011;
mem2[13133] = 10'b1111001011;
mem2[13134] = 10'b1111001011;
mem2[13135] = 10'b1111001011;
mem2[13136] = 10'b1111001011;
mem2[13137] = 10'b1111001100;
mem2[13138] = 10'b1111001100;
mem2[13139] = 10'b1111001100;
mem2[13140] = 10'b1111001100;
mem2[13141] = 10'b1111001100;
mem2[13142] = 10'b1111001100;
mem2[13143] = 10'b1111001100;
mem2[13144] = 10'b1111001100;
mem2[13145] = 10'b1111001100;
mem2[13146] = 10'b1111001100;
mem2[13147] = 10'b1111001100;
mem2[13148] = 10'b1111001100;
mem2[13149] = 10'b1111001100;
mem2[13150] = 10'b1111001100;
mem2[13151] = 10'b1111001100;
mem2[13152] = 10'b1111001100;
mem2[13153] = 10'b1111001100;
mem2[13154] = 10'b1111001100;
mem2[13155] = 10'b1111001100;
mem2[13156] = 10'b1111001100;
mem2[13157] = 10'b1111001100;
mem2[13158] = 10'b1111001100;
mem2[13159] = 10'b1111001101;
mem2[13160] = 10'b1111001101;
mem2[13161] = 10'b1111001101;
mem2[13162] = 10'b1111001101;
mem2[13163] = 10'b1111001101;
mem2[13164] = 10'b1111001101;
mem2[13165] = 10'b1111001101;
mem2[13166] = 10'b1111001101;
mem2[13167] = 10'b1111001101;
mem2[13168] = 10'b1111001101;
mem2[13169] = 10'b1111001101;
mem2[13170] = 10'b1111001101;
mem2[13171] = 10'b1111001101;
mem2[13172] = 10'b1111001101;
mem2[13173] = 10'b1111001101;
mem2[13174] = 10'b1111001101;
mem2[13175] = 10'b1111001101;
mem2[13176] = 10'b1111001101;
mem2[13177] = 10'b1111001101;
mem2[13178] = 10'b1111001101;
mem2[13179] = 10'b1111001101;
mem2[13180] = 10'b1111001101;
mem2[13181] = 10'b1111001110;
mem2[13182] = 10'b1111001110;
mem2[13183] = 10'b1111001110;
mem2[13184] = 10'b1111001110;
mem2[13185] = 10'b1111001110;
mem2[13186] = 10'b1111001110;
mem2[13187] = 10'b1111001110;
mem2[13188] = 10'b1111001110;
mem2[13189] = 10'b1111001110;
mem2[13190] = 10'b1111001110;
mem2[13191] = 10'b1111001110;
mem2[13192] = 10'b1111001110;
mem2[13193] = 10'b1111001110;
mem2[13194] = 10'b1111001110;
mem2[13195] = 10'b1111001110;
mem2[13196] = 10'b1111001110;
mem2[13197] = 10'b1111001110;
mem2[13198] = 10'b1111001110;
mem2[13199] = 10'b1111001110;
mem2[13200] = 10'b1111001110;
mem2[13201] = 10'b1111001110;
mem2[13202] = 10'b1111001110;
mem2[13203] = 10'b1111001111;
mem2[13204] = 10'b1111001111;
mem2[13205] = 10'b1111001111;
mem2[13206] = 10'b1111001111;
mem2[13207] = 10'b1111001111;
mem2[13208] = 10'b1111001111;
mem2[13209] = 10'b1111001111;
mem2[13210] = 10'b1111001111;
mem2[13211] = 10'b1111001111;
mem2[13212] = 10'b1111001111;
mem2[13213] = 10'b1111001111;
mem2[13214] = 10'b1111001111;
mem2[13215] = 10'b1111001111;
mem2[13216] = 10'b1111001111;
mem2[13217] = 10'b1111001111;
mem2[13218] = 10'b1111001111;
mem2[13219] = 10'b1111001111;
mem2[13220] = 10'b1111001111;
mem2[13221] = 10'b1111001111;
mem2[13222] = 10'b1111001111;
mem2[13223] = 10'b1111001111;
mem2[13224] = 10'b1111001111;
mem2[13225] = 10'b1111001111;
mem2[13226] = 10'b1111010000;
mem2[13227] = 10'b1111010000;
mem2[13228] = 10'b1111010000;
mem2[13229] = 10'b1111010000;
mem2[13230] = 10'b1111010000;
mem2[13231] = 10'b1111010000;
mem2[13232] = 10'b1111010000;
mem2[13233] = 10'b1111010000;
mem2[13234] = 10'b1111010000;
mem2[13235] = 10'b1111010000;
mem2[13236] = 10'b1111010000;
mem2[13237] = 10'b1111010000;
mem2[13238] = 10'b1111010000;
mem2[13239] = 10'b1111010000;
mem2[13240] = 10'b1111010000;
mem2[13241] = 10'b1111010000;
mem2[13242] = 10'b1111010000;
mem2[13243] = 10'b1111010000;
mem2[13244] = 10'b1111010000;
mem2[13245] = 10'b1111010000;
mem2[13246] = 10'b1111010000;
mem2[13247] = 10'b1111010000;
mem2[13248] = 10'b1111010000;
mem2[13249] = 10'b1111010001;
mem2[13250] = 10'b1111010001;
mem2[13251] = 10'b1111010001;
mem2[13252] = 10'b1111010001;
mem2[13253] = 10'b1111010001;
mem2[13254] = 10'b1111010001;
mem2[13255] = 10'b1111010001;
mem2[13256] = 10'b1111010001;
mem2[13257] = 10'b1111010001;
mem2[13258] = 10'b1111010001;
mem2[13259] = 10'b1111010001;
mem2[13260] = 10'b1111010001;
mem2[13261] = 10'b1111010001;
mem2[13262] = 10'b1111010001;
mem2[13263] = 10'b1111010001;
mem2[13264] = 10'b1111010001;
mem2[13265] = 10'b1111010001;
mem2[13266] = 10'b1111010001;
mem2[13267] = 10'b1111010001;
mem2[13268] = 10'b1111010001;
mem2[13269] = 10'b1111010001;
mem2[13270] = 10'b1111010001;
mem2[13271] = 10'b1111010010;
mem2[13272] = 10'b1111010010;
mem2[13273] = 10'b1111010010;
mem2[13274] = 10'b1111010010;
mem2[13275] = 10'b1111010010;
mem2[13276] = 10'b1111010010;
mem2[13277] = 10'b1111010010;
mem2[13278] = 10'b1111010010;
mem2[13279] = 10'b1111010010;
mem2[13280] = 10'b1111010010;
mem2[13281] = 10'b1111010010;
mem2[13282] = 10'b1111010010;
mem2[13283] = 10'b1111010010;
mem2[13284] = 10'b1111010010;
mem2[13285] = 10'b1111010010;
mem2[13286] = 10'b1111010010;
mem2[13287] = 10'b1111010010;
mem2[13288] = 10'b1111010010;
mem2[13289] = 10'b1111010010;
mem2[13290] = 10'b1111010010;
mem2[13291] = 10'b1111010010;
mem2[13292] = 10'b1111010010;
mem2[13293] = 10'b1111010010;
mem2[13294] = 10'b1111010010;
mem2[13295] = 10'b1111010011;
mem2[13296] = 10'b1111010011;
mem2[13297] = 10'b1111010011;
mem2[13298] = 10'b1111010011;
mem2[13299] = 10'b1111010011;
mem2[13300] = 10'b1111010011;
mem2[13301] = 10'b1111010011;
mem2[13302] = 10'b1111010011;
mem2[13303] = 10'b1111010011;
mem2[13304] = 10'b1111010011;
mem2[13305] = 10'b1111010011;
mem2[13306] = 10'b1111010011;
mem2[13307] = 10'b1111010011;
mem2[13308] = 10'b1111010011;
mem2[13309] = 10'b1111010011;
mem2[13310] = 10'b1111010011;
mem2[13311] = 10'b1111010011;
mem2[13312] = 10'b1111010011;
mem2[13313] = 10'b1111010011;
mem2[13314] = 10'b1111010011;
mem2[13315] = 10'b1111010011;
mem2[13316] = 10'b1111010011;
mem2[13317] = 10'b1111010011;
mem2[13318] = 10'b1111010100;
mem2[13319] = 10'b1111010100;
mem2[13320] = 10'b1111010100;
mem2[13321] = 10'b1111010100;
mem2[13322] = 10'b1111010100;
mem2[13323] = 10'b1111010100;
mem2[13324] = 10'b1111010100;
mem2[13325] = 10'b1111010100;
mem2[13326] = 10'b1111010100;
mem2[13327] = 10'b1111010100;
mem2[13328] = 10'b1111010100;
mem2[13329] = 10'b1111010100;
mem2[13330] = 10'b1111010100;
mem2[13331] = 10'b1111010100;
mem2[13332] = 10'b1111010100;
mem2[13333] = 10'b1111010100;
mem2[13334] = 10'b1111010100;
mem2[13335] = 10'b1111010100;
mem2[13336] = 10'b1111010100;
mem2[13337] = 10'b1111010100;
mem2[13338] = 10'b1111010100;
mem2[13339] = 10'b1111010100;
mem2[13340] = 10'b1111010100;
mem2[13341] = 10'b1111010100;
mem2[13342] = 10'b1111010101;
mem2[13343] = 10'b1111010101;
mem2[13344] = 10'b1111010101;
mem2[13345] = 10'b1111010101;
mem2[13346] = 10'b1111010101;
mem2[13347] = 10'b1111010101;
mem2[13348] = 10'b1111010101;
mem2[13349] = 10'b1111010101;
mem2[13350] = 10'b1111010101;
mem2[13351] = 10'b1111010101;
mem2[13352] = 10'b1111010101;
mem2[13353] = 10'b1111010101;
mem2[13354] = 10'b1111010101;
mem2[13355] = 10'b1111010101;
mem2[13356] = 10'b1111010101;
mem2[13357] = 10'b1111010101;
mem2[13358] = 10'b1111010101;
mem2[13359] = 10'b1111010101;
mem2[13360] = 10'b1111010101;
mem2[13361] = 10'b1111010101;
mem2[13362] = 10'b1111010101;
mem2[13363] = 10'b1111010101;
mem2[13364] = 10'b1111010101;
mem2[13365] = 10'b1111010101;
mem2[13366] = 10'b1111010110;
mem2[13367] = 10'b1111010110;
mem2[13368] = 10'b1111010110;
mem2[13369] = 10'b1111010110;
mem2[13370] = 10'b1111010110;
mem2[13371] = 10'b1111010110;
mem2[13372] = 10'b1111010110;
mem2[13373] = 10'b1111010110;
mem2[13374] = 10'b1111010110;
mem2[13375] = 10'b1111010110;
mem2[13376] = 10'b1111010110;
mem2[13377] = 10'b1111010110;
mem2[13378] = 10'b1111010110;
mem2[13379] = 10'b1111010110;
mem2[13380] = 10'b1111010110;
mem2[13381] = 10'b1111010110;
mem2[13382] = 10'b1111010110;
mem2[13383] = 10'b1111010110;
mem2[13384] = 10'b1111010110;
mem2[13385] = 10'b1111010110;
mem2[13386] = 10'b1111010110;
mem2[13387] = 10'b1111010110;
mem2[13388] = 10'b1111010110;
mem2[13389] = 10'b1111010110;
mem2[13390] = 10'b1111010111;
mem2[13391] = 10'b1111010111;
mem2[13392] = 10'b1111010111;
mem2[13393] = 10'b1111010111;
mem2[13394] = 10'b1111010111;
mem2[13395] = 10'b1111010111;
mem2[13396] = 10'b1111010111;
mem2[13397] = 10'b1111010111;
mem2[13398] = 10'b1111010111;
mem2[13399] = 10'b1111010111;
mem2[13400] = 10'b1111010111;
mem2[13401] = 10'b1111010111;
mem2[13402] = 10'b1111010111;
mem2[13403] = 10'b1111010111;
mem2[13404] = 10'b1111010111;
mem2[13405] = 10'b1111010111;
mem2[13406] = 10'b1111010111;
mem2[13407] = 10'b1111010111;
mem2[13408] = 10'b1111010111;
mem2[13409] = 10'b1111010111;
mem2[13410] = 10'b1111010111;
mem2[13411] = 10'b1111010111;
mem2[13412] = 10'b1111010111;
mem2[13413] = 10'b1111010111;
mem2[13414] = 10'b1111011000;
mem2[13415] = 10'b1111011000;
mem2[13416] = 10'b1111011000;
mem2[13417] = 10'b1111011000;
mem2[13418] = 10'b1111011000;
mem2[13419] = 10'b1111011000;
mem2[13420] = 10'b1111011000;
mem2[13421] = 10'b1111011000;
mem2[13422] = 10'b1111011000;
mem2[13423] = 10'b1111011000;
mem2[13424] = 10'b1111011000;
mem2[13425] = 10'b1111011000;
mem2[13426] = 10'b1111011000;
mem2[13427] = 10'b1111011000;
mem2[13428] = 10'b1111011000;
mem2[13429] = 10'b1111011000;
mem2[13430] = 10'b1111011000;
mem2[13431] = 10'b1111011000;
mem2[13432] = 10'b1111011000;
mem2[13433] = 10'b1111011000;
mem2[13434] = 10'b1111011000;
mem2[13435] = 10'b1111011000;
mem2[13436] = 10'b1111011000;
mem2[13437] = 10'b1111011000;
mem2[13438] = 10'b1111011000;
mem2[13439] = 10'b1111011001;
mem2[13440] = 10'b1111011001;
mem2[13441] = 10'b1111011001;
mem2[13442] = 10'b1111011001;
mem2[13443] = 10'b1111011001;
mem2[13444] = 10'b1111011001;
mem2[13445] = 10'b1111011001;
mem2[13446] = 10'b1111011001;
mem2[13447] = 10'b1111011001;
mem2[13448] = 10'b1111011001;
mem2[13449] = 10'b1111011001;
mem2[13450] = 10'b1111011001;
mem2[13451] = 10'b1111011001;
mem2[13452] = 10'b1111011001;
mem2[13453] = 10'b1111011001;
mem2[13454] = 10'b1111011001;
mem2[13455] = 10'b1111011001;
mem2[13456] = 10'b1111011001;
mem2[13457] = 10'b1111011001;
mem2[13458] = 10'b1111011001;
mem2[13459] = 10'b1111011001;
mem2[13460] = 10'b1111011001;
mem2[13461] = 10'b1111011001;
mem2[13462] = 10'b1111011001;
mem2[13463] = 10'b1111011001;
mem2[13464] = 10'b1111011010;
mem2[13465] = 10'b1111011010;
mem2[13466] = 10'b1111011010;
mem2[13467] = 10'b1111011010;
mem2[13468] = 10'b1111011010;
mem2[13469] = 10'b1111011010;
mem2[13470] = 10'b1111011010;
mem2[13471] = 10'b1111011010;
mem2[13472] = 10'b1111011010;
mem2[13473] = 10'b1111011010;
mem2[13474] = 10'b1111011010;
mem2[13475] = 10'b1111011010;
mem2[13476] = 10'b1111011010;
mem2[13477] = 10'b1111011010;
mem2[13478] = 10'b1111011010;
mem2[13479] = 10'b1111011010;
mem2[13480] = 10'b1111011010;
mem2[13481] = 10'b1111011010;
mem2[13482] = 10'b1111011010;
mem2[13483] = 10'b1111011010;
mem2[13484] = 10'b1111011010;
mem2[13485] = 10'b1111011010;
mem2[13486] = 10'b1111011010;
mem2[13487] = 10'b1111011010;
mem2[13488] = 10'b1111011010;
mem2[13489] = 10'b1111011010;
mem2[13490] = 10'b1111011011;
mem2[13491] = 10'b1111011011;
mem2[13492] = 10'b1111011011;
mem2[13493] = 10'b1111011011;
mem2[13494] = 10'b1111011011;
mem2[13495] = 10'b1111011011;
mem2[13496] = 10'b1111011011;
mem2[13497] = 10'b1111011011;
mem2[13498] = 10'b1111011011;
mem2[13499] = 10'b1111011011;
mem2[13500] = 10'b1111011011;
mem2[13501] = 10'b1111011011;
mem2[13502] = 10'b1111011011;
mem2[13503] = 10'b1111011011;
mem2[13504] = 10'b1111011011;
mem2[13505] = 10'b1111011011;
mem2[13506] = 10'b1111011011;
mem2[13507] = 10'b1111011011;
mem2[13508] = 10'b1111011011;
mem2[13509] = 10'b1111011011;
mem2[13510] = 10'b1111011011;
mem2[13511] = 10'b1111011011;
mem2[13512] = 10'b1111011011;
mem2[13513] = 10'b1111011011;
mem2[13514] = 10'b1111011011;
mem2[13515] = 10'b1111011100;
mem2[13516] = 10'b1111011100;
mem2[13517] = 10'b1111011100;
mem2[13518] = 10'b1111011100;
mem2[13519] = 10'b1111011100;
mem2[13520] = 10'b1111011100;
mem2[13521] = 10'b1111011100;
mem2[13522] = 10'b1111011100;
mem2[13523] = 10'b1111011100;
mem2[13524] = 10'b1111011100;
mem2[13525] = 10'b1111011100;
mem2[13526] = 10'b1111011100;
mem2[13527] = 10'b1111011100;
mem2[13528] = 10'b1111011100;
mem2[13529] = 10'b1111011100;
mem2[13530] = 10'b1111011100;
mem2[13531] = 10'b1111011100;
mem2[13532] = 10'b1111011100;
mem2[13533] = 10'b1111011100;
mem2[13534] = 10'b1111011100;
mem2[13535] = 10'b1111011100;
mem2[13536] = 10'b1111011100;
mem2[13537] = 10'b1111011100;
mem2[13538] = 10'b1111011100;
mem2[13539] = 10'b1111011100;
mem2[13540] = 10'b1111011100;
mem2[13541] = 10'b1111011100;
mem2[13542] = 10'b1111011101;
mem2[13543] = 10'b1111011101;
mem2[13544] = 10'b1111011101;
mem2[13545] = 10'b1111011101;
mem2[13546] = 10'b1111011101;
mem2[13547] = 10'b1111011101;
mem2[13548] = 10'b1111011101;
mem2[13549] = 10'b1111011101;
mem2[13550] = 10'b1111011101;
mem2[13551] = 10'b1111011101;
mem2[13552] = 10'b1111011101;
mem2[13553] = 10'b1111011101;
mem2[13554] = 10'b1111011101;
mem2[13555] = 10'b1111011101;
mem2[13556] = 10'b1111011101;
mem2[13557] = 10'b1111011101;
mem2[13558] = 10'b1111011101;
mem2[13559] = 10'b1111011101;
mem2[13560] = 10'b1111011101;
mem2[13561] = 10'b1111011101;
mem2[13562] = 10'b1111011101;
mem2[13563] = 10'b1111011101;
mem2[13564] = 10'b1111011101;
mem2[13565] = 10'b1111011101;
mem2[13566] = 10'b1111011101;
mem2[13567] = 10'b1111011101;
mem2[13568] = 10'b1111011110;
mem2[13569] = 10'b1111011110;
mem2[13570] = 10'b1111011110;
mem2[13571] = 10'b1111011110;
mem2[13572] = 10'b1111011110;
mem2[13573] = 10'b1111011110;
mem2[13574] = 10'b1111011110;
mem2[13575] = 10'b1111011110;
mem2[13576] = 10'b1111011110;
mem2[13577] = 10'b1111011110;
mem2[13578] = 10'b1111011110;
mem2[13579] = 10'b1111011110;
mem2[13580] = 10'b1111011110;
mem2[13581] = 10'b1111011110;
mem2[13582] = 10'b1111011110;
mem2[13583] = 10'b1111011110;
mem2[13584] = 10'b1111011110;
mem2[13585] = 10'b1111011110;
mem2[13586] = 10'b1111011110;
mem2[13587] = 10'b1111011110;
mem2[13588] = 10'b1111011110;
mem2[13589] = 10'b1111011110;
mem2[13590] = 10'b1111011110;
mem2[13591] = 10'b1111011110;
mem2[13592] = 10'b1111011110;
mem2[13593] = 10'b1111011110;
mem2[13594] = 10'b1111011110;
mem2[13595] = 10'b1111011111;
mem2[13596] = 10'b1111011111;
mem2[13597] = 10'b1111011111;
mem2[13598] = 10'b1111011111;
mem2[13599] = 10'b1111011111;
mem2[13600] = 10'b1111011111;
mem2[13601] = 10'b1111011111;
mem2[13602] = 10'b1111011111;
mem2[13603] = 10'b1111011111;
mem2[13604] = 10'b1111011111;
mem2[13605] = 10'b1111011111;
mem2[13606] = 10'b1111011111;
mem2[13607] = 10'b1111011111;
mem2[13608] = 10'b1111011111;
mem2[13609] = 10'b1111011111;
mem2[13610] = 10'b1111011111;
mem2[13611] = 10'b1111011111;
mem2[13612] = 10'b1111011111;
mem2[13613] = 10'b1111011111;
mem2[13614] = 10'b1111011111;
mem2[13615] = 10'b1111011111;
mem2[13616] = 10'b1111011111;
mem2[13617] = 10'b1111011111;
mem2[13618] = 10'b1111011111;
mem2[13619] = 10'b1111011111;
mem2[13620] = 10'b1111011111;
mem2[13621] = 10'b1111011111;
mem2[13622] = 10'b1111100000;
mem2[13623] = 10'b1111100000;
mem2[13624] = 10'b1111100000;
mem2[13625] = 10'b1111100000;
mem2[13626] = 10'b1111100000;
mem2[13627] = 10'b1111100000;
mem2[13628] = 10'b1111100000;
mem2[13629] = 10'b1111100000;
mem2[13630] = 10'b1111100000;
mem2[13631] = 10'b1111100000;
mem2[13632] = 10'b1111100000;
mem2[13633] = 10'b1111100000;
mem2[13634] = 10'b1111100000;
mem2[13635] = 10'b1111100000;
mem2[13636] = 10'b1111100000;
mem2[13637] = 10'b1111100000;
mem2[13638] = 10'b1111100000;
mem2[13639] = 10'b1111100000;
mem2[13640] = 10'b1111100000;
mem2[13641] = 10'b1111100000;
mem2[13642] = 10'b1111100000;
mem2[13643] = 10'b1111100000;
mem2[13644] = 10'b1111100000;
mem2[13645] = 10'b1111100000;
mem2[13646] = 10'b1111100000;
mem2[13647] = 10'b1111100000;
mem2[13648] = 10'b1111100000;
mem2[13649] = 10'b1111100000;
mem2[13650] = 10'b1111100001;
mem2[13651] = 10'b1111100001;
mem2[13652] = 10'b1111100001;
mem2[13653] = 10'b1111100001;
mem2[13654] = 10'b1111100001;
mem2[13655] = 10'b1111100001;
mem2[13656] = 10'b1111100001;
mem2[13657] = 10'b1111100001;
mem2[13658] = 10'b1111100001;
mem2[13659] = 10'b1111100001;
mem2[13660] = 10'b1111100001;
mem2[13661] = 10'b1111100001;
mem2[13662] = 10'b1111100001;
mem2[13663] = 10'b1111100001;
mem2[13664] = 10'b1111100001;
mem2[13665] = 10'b1111100001;
mem2[13666] = 10'b1111100001;
mem2[13667] = 10'b1111100001;
mem2[13668] = 10'b1111100001;
mem2[13669] = 10'b1111100001;
mem2[13670] = 10'b1111100001;
mem2[13671] = 10'b1111100001;
mem2[13672] = 10'b1111100001;
mem2[13673] = 10'b1111100001;
mem2[13674] = 10'b1111100001;
mem2[13675] = 10'b1111100001;
mem2[13676] = 10'b1111100001;
mem2[13677] = 10'b1111100001;
mem2[13678] = 10'b1111100010;
mem2[13679] = 10'b1111100010;
mem2[13680] = 10'b1111100010;
mem2[13681] = 10'b1111100010;
mem2[13682] = 10'b1111100010;
mem2[13683] = 10'b1111100010;
mem2[13684] = 10'b1111100010;
mem2[13685] = 10'b1111100010;
mem2[13686] = 10'b1111100010;
mem2[13687] = 10'b1111100010;
mem2[13688] = 10'b1111100010;
mem2[13689] = 10'b1111100010;
mem2[13690] = 10'b1111100010;
mem2[13691] = 10'b1111100010;
mem2[13692] = 10'b1111100010;
mem2[13693] = 10'b1111100010;
mem2[13694] = 10'b1111100010;
mem2[13695] = 10'b1111100010;
mem2[13696] = 10'b1111100010;
mem2[13697] = 10'b1111100010;
mem2[13698] = 10'b1111100010;
mem2[13699] = 10'b1111100010;
mem2[13700] = 10'b1111100010;
mem2[13701] = 10'b1111100010;
mem2[13702] = 10'b1111100010;
mem2[13703] = 10'b1111100010;
mem2[13704] = 10'b1111100010;
mem2[13705] = 10'b1111100010;
mem2[13706] = 10'b1111100011;
mem2[13707] = 10'b1111100011;
mem2[13708] = 10'b1111100011;
mem2[13709] = 10'b1111100011;
mem2[13710] = 10'b1111100011;
mem2[13711] = 10'b1111100011;
mem2[13712] = 10'b1111100011;
mem2[13713] = 10'b1111100011;
mem2[13714] = 10'b1111100011;
mem2[13715] = 10'b1111100011;
mem2[13716] = 10'b1111100011;
mem2[13717] = 10'b1111100011;
mem2[13718] = 10'b1111100011;
mem2[13719] = 10'b1111100011;
mem2[13720] = 10'b1111100011;
mem2[13721] = 10'b1111100011;
mem2[13722] = 10'b1111100011;
mem2[13723] = 10'b1111100011;
mem2[13724] = 10'b1111100011;
mem2[13725] = 10'b1111100011;
mem2[13726] = 10'b1111100011;
mem2[13727] = 10'b1111100011;
mem2[13728] = 10'b1111100011;
mem2[13729] = 10'b1111100011;
mem2[13730] = 10'b1111100011;
mem2[13731] = 10'b1111100011;
mem2[13732] = 10'b1111100011;
mem2[13733] = 10'b1111100011;
mem2[13734] = 10'b1111100011;
mem2[13735] = 10'b1111100100;
mem2[13736] = 10'b1111100100;
mem2[13737] = 10'b1111100100;
mem2[13738] = 10'b1111100100;
mem2[13739] = 10'b1111100100;
mem2[13740] = 10'b1111100100;
mem2[13741] = 10'b1111100100;
mem2[13742] = 10'b1111100100;
mem2[13743] = 10'b1111100100;
mem2[13744] = 10'b1111100100;
mem2[13745] = 10'b1111100100;
mem2[13746] = 10'b1111100100;
mem2[13747] = 10'b1111100100;
mem2[13748] = 10'b1111100100;
mem2[13749] = 10'b1111100100;
mem2[13750] = 10'b1111100100;
mem2[13751] = 10'b1111100100;
mem2[13752] = 10'b1111100100;
mem2[13753] = 10'b1111100100;
mem2[13754] = 10'b1111100100;
mem2[13755] = 10'b1111100100;
mem2[13756] = 10'b1111100100;
mem2[13757] = 10'b1111100100;
mem2[13758] = 10'b1111100100;
mem2[13759] = 10'b1111100100;
mem2[13760] = 10'b1111100100;
mem2[13761] = 10'b1111100100;
mem2[13762] = 10'b1111100100;
mem2[13763] = 10'b1111100100;
mem2[13764] = 10'b1111100100;
mem2[13765] = 10'b1111100101;
mem2[13766] = 10'b1111100101;
mem2[13767] = 10'b1111100101;
mem2[13768] = 10'b1111100101;
mem2[13769] = 10'b1111100101;
mem2[13770] = 10'b1111100101;
mem2[13771] = 10'b1111100101;
mem2[13772] = 10'b1111100101;
mem2[13773] = 10'b1111100101;
mem2[13774] = 10'b1111100101;
mem2[13775] = 10'b1111100101;
mem2[13776] = 10'b1111100101;
mem2[13777] = 10'b1111100101;
mem2[13778] = 10'b1111100101;
mem2[13779] = 10'b1111100101;
mem2[13780] = 10'b1111100101;
mem2[13781] = 10'b1111100101;
mem2[13782] = 10'b1111100101;
mem2[13783] = 10'b1111100101;
mem2[13784] = 10'b1111100101;
mem2[13785] = 10'b1111100101;
mem2[13786] = 10'b1111100101;
mem2[13787] = 10'b1111100101;
mem2[13788] = 10'b1111100101;
mem2[13789] = 10'b1111100101;
mem2[13790] = 10'b1111100101;
mem2[13791] = 10'b1111100101;
mem2[13792] = 10'b1111100101;
mem2[13793] = 10'b1111100101;
mem2[13794] = 10'b1111100101;
mem2[13795] = 10'b1111100110;
mem2[13796] = 10'b1111100110;
mem2[13797] = 10'b1111100110;
mem2[13798] = 10'b1111100110;
mem2[13799] = 10'b1111100110;
mem2[13800] = 10'b1111100110;
mem2[13801] = 10'b1111100110;
mem2[13802] = 10'b1111100110;
mem2[13803] = 10'b1111100110;
mem2[13804] = 10'b1111100110;
mem2[13805] = 10'b1111100110;
mem2[13806] = 10'b1111100110;
mem2[13807] = 10'b1111100110;
mem2[13808] = 10'b1111100110;
mem2[13809] = 10'b1111100110;
mem2[13810] = 10'b1111100110;
mem2[13811] = 10'b1111100110;
mem2[13812] = 10'b1111100110;
mem2[13813] = 10'b1111100110;
mem2[13814] = 10'b1111100110;
mem2[13815] = 10'b1111100110;
mem2[13816] = 10'b1111100110;
mem2[13817] = 10'b1111100110;
mem2[13818] = 10'b1111100110;
mem2[13819] = 10'b1111100110;
mem2[13820] = 10'b1111100110;
mem2[13821] = 10'b1111100110;
mem2[13822] = 10'b1111100110;
mem2[13823] = 10'b1111100110;
mem2[13824] = 10'b1111100110;
mem2[13825] = 10'b1111100110;
mem2[13826] = 10'b1111100111;
mem2[13827] = 10'b1111100111;
mem2[13828] = 10'b1111100111;
mem2[13829] = 10'b1111100111;
mem2[13830] = 10'b1111100111;
mem2[13831] = 10'b1111100111;
mem2[13832] = 10'b1111100111;
mem2[13833] = 10'b1111100111;
mem2[13834] = 10'b1111100111;
mem2[13835] = 10'b1111100111;
mem2[13836] = 10'b1111100111;
mem2[13837] = 10'b1111100111;
mem2[13838] = 10'b1111100111;
mem2[13839] = 10'b1111100111;
mem2[13840] = 10'b1111100111;
mem2[13841] = 10'b1111100111;
mem2[13842] = 10'b1111100111;
mem2[13843] = 10'b1111100111;
mem2[13844] = 10'b1111100111;
mem2[13845] = 10'b1111100111;
mem2[13846] = 10'b1111100111;
mem2[13847] = 10'b1111100111;
mem2[13848] = 10'b1111100111;
mem2[13849] = 10'b1111100111;
mem2[13850] = 10'b1111100111;
mem2[13851] = 10'b1111100111;
mem2[13852] = 10'b1111100111;
mem2[13853] = 10'b1111100111;
mem2[13854] = 10'b1111100111;
mem2[13855] = 10'b1111100111;
mem2[13856] = 10'b1111100111;
mem2[13857] = 10'b1111101000;
mem2[13858] = 10'b1111101000;
mem2[13859] = 10'b1111101000;
mem2[13860] = 10'b1111101000;
mem2[13861] = 10'b1111101000;
mem2[13862] = 10'b1111101000;
mem2[13863] = 10'b1111101000;
mem2[13864] = 10'b1111101000;
mem2[13865] = 10'b1111101000;
mem2[13866] = 10'b1111101000;
mem2[13867] = 10'b1111101000;
mem2[13868] = 10'b1111101000;
mem2[13869] = 10'b1111101000;
mem2[13870] = 10'b1111101000;
mem2[13871] = 10'b1111101000;
mem2[13872] = 10'b1111101000;
mem2[13873] = 10'b1111101000;
mem2[13874] = 10'b1111101000;
mem2[13875] = 10'b1111101000;
mem2[13876] = 10'b1111101000;
mem2[13877] = 10'b1111101000;
mem2[13878] = 10'b1111101000;
mem2[13879] = 10'b1111101000;
mem2[13880] = 10'b1111101000;
mem2[13881] = 10'b1111101000;
mem2[13882] = 10'b1111101000;
mem2[13883] = 10'b1111101000;
mem2[13884] = 10'b1111101000;
mem2[13885] = 10'b1111101000;
mem2[13886] = 10'b1111101000;
mem2[13887] = 10'b1111101000;
mem2[13888] = 10'b1111101000;
mem2[13889] = 10'b1111101001;
mem2[13890] = 10'b1111101001;
mem2[13891] = 10'b1111101001;
mem2[13892] = 10'b1111101001;
mem2[13893] = 10'b1111101001;
mem2[13894] = 10'b1111101001;
mem2[13895] = 10'b1111101001;
mem2[13896] = 10'b1111101001;
mem2[13897] = 10'b1111101001;
mem2[13898] = 10'b1111101001;
mem2[13899] = 10'b1111101001;
mem2[13900] = 10'b1111101001;
mem2[13901] = 10'b1111101001;
mem2[13902] = 10'b1111101001;
mem2[13903] = 10'b1111101001;
mem2[13904] = 10'b1111101001;
mem2[13905] = 10'b1111101001;
mem2[13906] = 10'b1111101001;
mem2[13907] = 10'b1111101001;
mem2[13908] = 10'b1111101001;
mem2[13909] = 10'b1111101001;
mem2[13910] = 10'b1111101001;
mem2[13911] = 10'b1111101001;
mem2[13912] = 10'b1111101001;
mem2[13913] = 10'b1111101001;
mem2[13914] = 10'b1111101001;
mem2[13915] = 10'b1111101001;
mem2[13916] = 10'b1111101001;
mem2[13917] = 10'b1111101001;
mem2[13918] = 10'b1111101001;
mem2[13919] = 10'b1111101001;
mem2[13920] = 10'b1111101001;
mem2[13921] = 10'b1111101010;
mem2[13922] = 10'b1111101010;
mem2[13923] = 10'b1111101010;
mem2[13924] = 10'b1111101010;
mem2[13925] = 10'b1111101010;
mem2[13926] = 10'b1111101010;
mem2[13927] = 10'b1111101010;
mem2[13928] = 10'b1111101010;
mem2[13929] = 10'b1111101010;
mem2[13930] = 10'b1111101010;
mem2[13931] = 10'b1111101010;
mem2[13932] = 10'b1111101010;
mem2[13933] = 10'b1111101010;
mem2[13934] = 10'b1111101010;
mem2[13935] = 10'b1111101010;
mem2[13936] = 10'b1111101010;
mem2[13937] = 10'b1111101010;
mem2[13938] = 10'b1111101010;
mem2[13939] = 10'b1111101010;
mem2[13940] = 10'b1111101010;
mem2[13941] = 10'b1111101010;
mem2[13942] = 10'b1111101010;
mem2[13943] = 10'b1111101010;
mem2[13944] = 10'b1111101010;
mem2[13945] = 10'b1111101010;
mem2[13946] = 10'b1111101010;
mem2[13947] = 10'b1111101010;
mem2[13948] = 10'b1111101010;
mem2[13949] = 10'b1111101010;
mem2[13950] = 10'b1111101010;
mem2[13951] = 10'b1111101010;
mem2[13952] = 10'b1111101010;
mem2[13953] = 10'b1111101010;
mem2[13954] = 10'b1111101010;
mem2[13955] = 10'b1111101011;
mem2[13956] = 10'b1111101011;
mem2[13957] = 10'b1111101011;
mem2[13958] = 10'b1111101011;
mem2[13959] = 10'b1111101011;
mem2[13960] = 10'b1111101011;
mem2[13961] = 10'b1111101011;
mem2[13962] = 10'b1111101011;
mem2[13963] = 10'b1111101011;
mem2[13964] = 10'b1111101011;
mem2[13965] = 10'b1111101011;
mem2[13966] = 10'b1111101011;
mem2[13967] = 10'b1111101011;
mem2[13968] = 10'b1111101011;
mem2[13969] = 10'b1111101011;
mem2[13970] = 10'b1111101011;
mem2[13971] = 10'b1111101011;
mem2[13972] = 10'b1111101011;
mem2[13973] = 10'b1111101011;
mem2[13974] = 10'b1111101011;
mem2[13975] = 10'b1111101011;
mem2[13976] = 10'b1111101011;
mem2[13977] = 10'b1111101011;
mem2[13978] = 10'b1111101011;
mem2[13979] = 10'b1111101011;
mem2[13980] = 10'b1111101011;
mem2[13981] = 10'b1111101011;
mem2[13982] = 10'b1111101011;
mem2[13983] = 10'b1111101011;
mem2[13984] = 10'b1111101011;
mem2[13985] = 10'b1111101011;
mem2[13986] = 10'b1111101011;
mem2[13987] = 10'b1111101011;
mem2[13988] = 10'b1111101011;
mem2[13989] = 10'b1111101100;
mem2[13990] = 10'b1111101100;
mem2[13991] = 10'b1111101100;
mem2[13992] = 10'b1111101100;
mem2[13993] = 10'b1111101100;
mem2[13994] = 10'b1111101100;
mem2[13995] = 10'b1111101100;
mem2[13996] = 10'b1111101100;
mem2[13997] = 10'b1111101100;
mem2[13998] = 10'b1111101100;
mem2[13999] = 10'b1111101100;
mem2[14000] = 10'b1111101100;
mem2[14001] = 10'b1111101100;
mem2[14002] = 10'b1111101100;
mem2[14003] = 10'b1111101100;
mem2[14004] = 10'b1111101100;
mem2[14005] = 10'b1111101100;
mem2[14006] = 10'b1111101100;
mem2[14007] = 10'b1111101100;
mem2[14008] = 10'b1111101100;
mem2[14009] = 10'b1111101100;
mem2[14010] = 10'b1111101100;
mem2[14011] = 10'b1111101100;
mem2[14012] = 10'b1111101100;
mem2[14013] = 10'b1111101100;
mem2[14014] = 10'b1111101100;
mem2[14015] = 10'b1111101100;
mem2[14016] = 10'b1111101100;
mem2[14017] = 10'b1111101100;
mem2[14018] = 10'b1111101100;
mem2[14019] = 10'b1111101100;
mem2[14020] = 10'b1111101100;
mem2[14021] = 10'b1111101100;
mem2[14022] = 10'b1111101100;
mem2[14023] = 10'b1111101100;
mem2[14024] = 10'b1111101101;
mem2[14025] = 10'b1111101101;
mem2[14026] = 10'b1111101101;
mem2[14027] = 10'b1111101101;
mem2[14028] = 10'b1111101101;
mem2[14029] = 10'b1111101101;
mem2[14030] = 10'b1111101101;
mem2[14031] = 10'b1111101101;
mem2[14032] = 10'b1111101101;
mem2[14033] = 10'b1111101101;
mem2[14034] = 10'b1111101101;
mem2[14035] = 10'b1111101101;
mem2[14036] = 10'b1111101101;
mem2[14037] = 10'b1111101101;
mem2[14038] = 10'b1111101101;
mem2[14039] = 10'b1111101101;
mem2[14040] = 10'b1111101101;
mem2[14041] = 10'b1111101101;
mem2[14042] = 10'b1111101101;
mem2[14043] = 10'b1111101101;
mem2[14044] = 10'b1111101101;
mem2[14045] = 10'b1111101101;
mem2[14046] = 10'b1111101101;
mem2[14047] = 10'b1111101101;
mem2[14048] = 10'b1111101101;
mem2[14049] = 10'b1111101101;
mem2[14050] = 10'b1111101101;
mem2[14051] = 10'b1111101101;
mem2[14052] = 10'b1111101101;
mem2[14053] = 10'b1111101101;
mem2[14054] = 10'b1111101101;
mem2[14055] = 10'b1111101101;
mem2[14056] = 10'b1111101101;
mem2[14057] = 10'b1111101101;
mem2[14058] = 10'b1111101101;
mem2[14059] = 10'b1111101101;
mem2[14060] = 10'b1111101110;
mem2[14061] = 10'b1111101110;
mem2[14062] = 10'b1111101110;
mem2[14063] = 10'b1111101110;
mem2[14064] = 10'b1111101110;
mem2[14065] = 10'b1111101110;
mem2[14066] = 10'b1111101110;
mem2[14067] = 10'b1111101110;
mem2[14068] = 10'b1111101110;
mem2[14069] = 10'b1111101110;
mem2[14070] = 10'b1111101110;
mem2[14071] = 10'b1111101110;
mem2[14072] = 10'b1111101110;
mem2[14073] = 10'b1111101110;
mem2[14074] = 10'b1111101110;
mem2[14075] = 10'b1111101110;
mem2[14076] = 10'b1111101110;
mem2[14077] = 10'b1111101110;
mem2[14078] = 10'b1111101110;
mem2[14079] = 10'b1111101110;
mem2[14080] = 10'b1111101110;
mem2[14081] = 10'b1111101110;
mem2[14082] = 10'b1111101110;
mem2[14083] = 10'b1111101110;
mem2[14084] = 10'b1111101110;
mem2[14085] = 10'b1111101110;
mem2[14086] = 10'b1111101110;
mem2[14087] = 10'b1111101110;
mem2[14088] = 10'b1111101110;
mem2[14089] = 10'b1111101110;
mem2[14090] = 10'b1111101110;
mem2[14091] = 10'b1111101110;
mem2[14092] = 10'b1111101110;
mem2[14093] = 10'b1111101110;
mem2[14094] = 10'b1111101110;
mem2[14095] = 10'b1111101110;
mem2[14096] = 10'b1111101111;
mem2[14097] = 10'b1111101111;
mem2[14098] = 10'b1111101111;
mem2[14099] = 10'b1111101111;
mem2[14100] = 10'b1111101111;
mem2[14101] = 10'b1111101111;
mem2[14102] = 10'b1111101111;
mem2[14103] = 10'b1111101111;
mem2[14104] = 10'b1111101111;
mem2[14105] = 10'b1111101111;
mem2[14106] = 10'b1111101111;
mem2[14107] = 10'b1111101111;
mem2[14108] = 10'b1111101111;
mem2[14109] = 10'b1111101111;
mem2[14110] = 10'b1111101111;
mem2[14111] = 10'b1111101111;
mem2[14112] = 10'b1111101111;
mem2[14113] = 10'b1111101111;
mem2[14114] = 10'b1111101111;
mem2[14115] = 10'b1111101111;
mem2[14116] = 10'b1111101111;
mem2[14117] = 10'b1111101111;
mem2[14118] = 10'b1111101111;
mem2[14119] = 10'b1111101111;
mem2[14120] = 10'b1111101111;
mem2[14121] = 10'b1111101111;
mem2[14122] = 10'b1111101111;
mem2[14123] = 10'b1111101111;
mem2[14124] = 10'b1111101111;
mem2[14125] = 10'b1111101111;
mem2[14126] = 10'b1111101111;
mem2[14127] = 10'b1111101111;
mem2[14128] = 10'b1111101111;
mem2[14129] = 10'b1111101111;
mem2[14130] = 10'b1111101111;
mem2[14131] = 10'b1111101111;
mem2[14132] = 10'b1111101111;
mem2[14133] = 10'b1111101111;
mem2[14134] = 10'b1111110000;
mem2[14135] = 10'b1111110000;
mem2[14136] = 10'b1111110000;
mem2[14137] = 10'b1111110000;
mem2[14138] = 10'b1111110000;
mem2[14139] = 10'b1111110000;
mem2[14140] = 10'b1111110000;
mem2[14141] = 10'b1111110000;
mem2[14142] = 10'b1111110000;
mem2[14143] = 10'b1111110000;
mem2[14144] = 10'b1111110000;
mem2[14145] = 10'b1111110000;
mem2[14146] = 10'b1111110000;
mem2[14147] = 10'b1111110000;
mem2[14148] = 10'b1111110000;
mem2[14149] = 10'b1111110000;
mem2[14150] = 10'b1111110000;
mem2[14151] = 10'b1111110000;
mem2[14152] = 10'b1111110000;
mem2[14153] = 10'b1111110000;
mem2[14154] = 10'b1111110000;
mem2[14155] = 10'b1111110000;
mem2[14156] = 10'b1111110000;
mem2[14157] = 10'b1111110000;
mem2[14158] = 10'b1111110000;
mem2[14159] = 10'b1111110000;
mem2[14160] = 10'b1111110000;
mem2[14161] = 10'b1111110000;
mem2[14162] = 10'b1111110000;
mem2[14163] = 10'b1111110000;
mem2[14164] = 10'b1111110000;
mem2[14165] = 10'b1111110000;
mem2[14166] = 10'b1111110000;
mem2[14167] = 10'b1111110000;
mem2[14168] = 10'b1111110000;
mem2[14169] = 10'b1111110000;
mem2[14170] = 10'b1111110000;
mem2[14171] = 10'b1111110000;
mem2[14172] = 10'b1111110000;
mem2[14173] = 10'b1111110001;
mem2[14174] = 10'b1111110001;
mem2[14175] = 10'b1111110001;
mem2[14176] = 10'b1111110001;
mem2[14177] = 10'b1111110001;
mem2[14178] = 10'b1111110001;
mem2[14179] = 10'b1111110001;
mem2[14180] = 10'b1111110001;
mem2[14181] = 10'b1111110001;
mem2[14182] = 10'b1111110001;
mem2[14183] = 10'b1111110001;
mem2[14184] = 10'b1111110001;
mem2[14185] = 10'b1111110001;
mem2[14186] = 10'b1111110001;
mem2[14187] = 10'b1111110001;
mem2[14188] = 10'b1111110001;
mem2[14189] = 10'b1111110001;
mem2[14190] = 10'b1111110001;
mem2[14191] = 10'b1111110001;
mem2[14192] = 10'b1111110001;
mem2[14193] = 10'b1111110001;
mem2[14194] = 10'b1111110001;
mem2[14195] = 10'b1111110001;
mem2[14196] = 10'b1111110001;
mem2[14197] = 10'b1111110001;
mem2[14198] = 10'b1111110001;
mem2[14199] = 10'b1111110001;
mem2[14200] = 10'b1111110001;
mem2[14201] = 10'b1111110001;
mem2[14202] = 10'b1111110001;
mem2[14203] = 10'b1111110001;
mem2[14204] = 10'b1111110001;
mem2[14205] = 10'b1111110001;
mem2[14206] = 10'b1111110001;
mem2[14207] = 10'b1111110001;
mem2[14208] = 10'b1111110001;
mem2[14209] = 10'b1111110001;
mem2[14210] = 10'b1111110001;
mem2[14211] = 10'b1111110001;
mem2[14212] = 10'b1111110001;
mem2[14213] = 10'b1111110001;
mem2[14214] = 10'b1111110010;
mem2[14215] = 10'b1111110010;
mem2[14216] = 10'b1111110010;
mem2[14217] = 10'b1111110010;
mem2[14218] = 10'b1111110010;
mem2[14219] = 10'b1111110010;
mem2[14220] = 10'b1111110010;
mem2[14221] = 10'b1111110010;
mem2[14222] = 10'b1111110010;
mem2[14223] = 10'b1111110010;
mem2[14224] = 10'b1111110010;
mem2[14225] = 10'b1111110010;
mem2[14226] = 10'b1111110010;
mem2[14227] = 10'b1111110010;
mem2[14228] = 10'b1111110010;
mem2[14229] = 10'b1111110010;
mem2[14230] = 10'b1111110010;
mem2[14231] = 10'b1111110010;
mem2[14232] = 10'b1111110010;
mem2[14233] = 10'b1111110010;
mem2[14234] = 10'b1111110010;
mem2[14235] = 10'b1111110010;
mem2[14236] = 10'b1111110010;
mem2[14237] = 10'b1111110010;
mem2[14238] = 10'b1111110010;
mem2[14239] = 10'b1111110010;
mem2[14240] = 10'b1111110010;
mem2[14241] = 10'b1111110010;
mem2[14242] = 10'b1111110010;
mem2[14243] = 10'b1111110010;
mem2[14244] = 10'b1111110010;
mem2[14245] = 10'b1111110010;
mem2[14246] = 10'b1111110010;
mem2[14247] = 10'b1111110010;
mem2[14248] = 10'b1111110010;
mem2[14249] = 10'b1111110010;
mem2[14250] = 10'b1111110010;
mem2[14251] = 10'b1111110010;
mem2[14252] = 10'b1111110010;
mem2[14253] = 10'b1111110010;
mem2[14254] = 10'b1111110010;
mem2[14255] = 10'b1111110010;
mem2[14256] = 10'b1111110011;
mem2[14257] = 10'b1111110011;
mem2[14258] = 10'b1111110011;
mem2[14259] = 10'b1111110011;
mem2[14260] = 10'b1111110011;
mem2[14261] = 10'b1111110011;
mem2[14262] = 10'b1111110011;
mem2[14263] = 10'b1111110011;
mem2[14264] = 10'b1111110011;
mem2[14265] = 10'b1111110011;
mem2[14266] = 10'b1111110011;
mem2[14267] = 10'b1111110011;
mem2[14268] = 10'b1111110011;
mem2[14269] = 10'b1111110011;
mem2[14270] = 10'b1111110011;
mem2[14271] = 10'b1111110011;
mem2[14272] = 10'b1111110011;
mem2[14273] = 10'b1111110011;
mem2[14274] = 10'b1111110011;
mem2[14275] = 10'b1111110011;
mem2[14276] = 10'b1111110011;
mem2[14277] = 10'b1111110011;
mem2[14278] = 10'b1111110011;
mem2[14279] = 10'b1111110011;
mem2[14280] = 10'b1111110011;
mem2[14281] = 10'b1111110011;
mem2[14282] = 10'b1111110011;
mem2[14283] = 10'b1111110011;
mem2[14284] = 10'b1111110011;
mem2[14285] = 10'b1111110011;
mem2[14286] = 10'b1111110011;
mem2[14287] = 10'b1111110011;
mem2[14288] = 10'b1111110011;
mem2[14289] = 10'b1111110011;
mem2[14290] = 10'b1111110011;
mem2[14291] = 10'b1111110011;
mem2[14292] = 10'b1111110011;
mem2[14293] = 10'b1111110011;
mem2[14294] = 10'b1111110011;
mem2[14295] = 10'b1111110011;
mem2[14296] = 10'b1111110011;
mem2[14297] = 10'b1111110011;
mem2[14298] = 10'b1111110011;
mem2[14299] = 10'b1111110100;
mem2[14300] = 10'b1111110100;
mem2[14301] = 10'b1111110100;
mem2[14302] = 10'b1111110100;
mem2[14303] = 10'b1111110100;
mem2[14304] = 10'b1111110100;
mem2[14305] = 10'b1111110100;
mem2[14306] = 10'b1111110100;
mem2[14307] = 10'b1111110100;
mem2[14308] = 10'b1111110100;
mem2[14309] = 10'b1111110100;
mem2[14310] = 10'b1111110100;
mem2[14311] = 10'b1111110100;
mem2[14312] = 10'b1111110100;
mem2[14313] = 10'b1111110100;
mem2[14314] = 10'b1111110100;
mem2[14315] = 10'b1111110100;
mem2[14316] = 10'b1111110100;
mem2[14317] = 10'b1111110100;
mem2[14318] = 10'b1111110100;
mem2[14319] = 10'b1111110100;
mem2[14320] = 10'b1111110100;
mem2[14321] = 10'b1111110100;
mem2[14322] = 10'b1111110100;
mem2[14323] = 10'b1111110100;
mem2[14324] = 10'b1111110100;
mem2[14325] = 10'b1111110100;
mem2[14326] = 10'b1111110100;
mem2[14327] = 10'b1111110100;
mem2[14328] = 10'b1111110100;
mem2[14329] = 10'b1111110100;
mem2[14330] = 10'b1111110100;
mem2[14331] = 10'b1111110100;
mem2[14332] = 10'b1111110100;
mem2[14333] = 10'b1111110100;
mem2[14334] = 10'b1111110100;
mem2[14335] = 10'b1111110100;
mem2[14336] = 10'b1111110100;
mem2[14337] = 10'b1111110100;
mem2[14338] = 10'b1111110100;
mem2[14339] = 10'b1111110100;
mem2[14340] = 10'b1111110100;
mem2[14341] = 10'b1111110100;
mem2[14342] = 10'b1111110100;
mem2[14343] = 10'b1111110100;
mem2[14344] = 10'b1111110101;
mem2[14345] = 10'b1111110101;
mem2[14346] = 10'b1111110101;
mem2[14347] = 10'b1111110101;
mem2[14348] = 10'b1111110101;
mem2[14349] = 10'b1111110101;
mem2[14350] = 10'b1111110101;
mem2[14351] = 10'b1111110101;
mem2[14352] = 10'b1111110101;
mem2[14353] = 10'b1111110101;
mem2[14354] = 10'b1111110101;
mem2[14355] = 10'b1111110101;
mem2[14356] = 10'b1111110101;
mem2[14357] = 10'b1111110101;
mem2[14358] = 10'b1111110101;
mem2[14359] = 10'b1111110101;
mem2[14360] = 10'b1111110101;
mem2[14361] = 10'b1111110101;
mem2[14362] = 10'b1111110101;
mem2[14363] = 10'b1111110101;
mem2[14364] = 10'b1111110101;
mem2[14365] = 10'b1111110101;
mem2[14366] = 10'b1111110101;
mem2[14367] = 10'b1111110101;
mem2[14368] = 10'b1111110101;
mem2[14369] = 10'b1111110101;
mem2[14370] = 10'b1111110101;
mem2[14371] = 10'b1111110101;
mem2[14372] = 10'b1111110101;
mem2[14373] = 10'b1111110101;
mem2[14374] = 10'b1111110101;
mem2[14375] = 10'b1111110101;
mem2[14376] = 10'b1111110101;
mem2[14377] = 10'b1111110101;
mem2[14378] = 10'b1111110101;
mem2[14379] = 10'b1111110101;
mem2[14380] = 10'b1111110101;
mem2[14381] = 10'b1111110101;
mem2[14382] = 10'b1111110101;
mem2[14383] = 10'b1111110101;
mem2[14384] = 10'b1111110101;
mem2[14385] = 10'b1111110101;
mem2[14386] = 10'b1111110101;
mem2[14387] = 10'b1111110101;
mem2[14388] = 10'b1111110101;
mem2[14389] = 10'b1111110101;
mem2[14390] = 10'b1111110101;
mem2[14391] = 10'b1111110101;
mem2[14392] = 10'b1111110110;
mem2[14393] = 10'b1111110110;
mem2[14394] = 10'b1111110110;
mem2[14395] = 10'b1111110110;
mem2[14396] = 10'b1111110110;
mem2[14397] = 10'b1111110110;
mem2[14398] = 10'b1111110110;
mem2[14399] = 10'b1111110110;
mem2[14400] = 10'b1111110110;
mem2[14401] = 10'b1111110110;
mem2[14402] = 10'b1111110110;
mem2[14403] = 10'b1111110110;
mem2[14404] = 10'b1111110110;
mem2[14405] = 10'b1111110110;
mem2[14406] = 10'b1111110110;
mem2[14407] = 10'b1111110110;
mem2[14408] = 10'b1111110110;
mem2[14409] = 10'b1111110110;
mem2[14410] = 10'b1111110110;
mem2[14411] = 10'b1111110110;
mem2[14412] = 10'b1111110110;
mem2[14413] = 10'b1111110110;
mem2[14414] = 10'b1111110110;
mem2[14415] = 10'b1111110110;
mem2[14416] = 10'b1111110110;
mem2[14417] = 10'b1111110110;
mem2[14418] = 10'b1111110110;
mem2[14419] = 10'b1111110110;
mem2[14420] = 10'b1111110110;
mem2[14421] = 10'b1111110110;
mem2[14422] = 10'b1111110110;
mem2[14423] = 10'b1111110110;
mem2[14424] = 10'b1111110110;
mem2[14425] = 10'b1111110110;
mem2[14426] = 10'b1111110110;
mem2[14427] = 10'b1111110110;
mem2[14428] = 10'b1111110110;
mem2[14429] = 10'b1111110110;
mem2[14430] = 10'b1111110110;
mem2[14431] = 10'b1111110110;
mem2[14432] = 10'b1111110110;
mem2[14433] = 10'b1111110110;
mem2[14434] = 10'b1111110110;
mem2[14435] = 10'b1111110110;
mem2[14436] = 10'b1111110110;
mem2[14437] = 10'b1111110110;
mem2[14438] = 10'b1111110110;
mem2[14439] = 10'b1111110110;
mem2[14440] = 10'b1111110110;
mem2[14441] = 10'b1111110110;
mem2[14442] = 10'b1111110111;
mem2[14443] = 10'b1111110111;
mem2[14444] = 10'b1111110111;
mem2[14445] = 10'b1111110111;
mem2[14446] = 10'b1111110111;
mem2[14447] = 10'b1111110111;
mem2[14448] = 10'b1111110111;
mem2[14449] = 10'b1111110111;
mem2[14450] = 10'b1111110111;
mem2[14451] = 10'b1111110111;
mem2[14452] = 10'b1111110111;
mem2[14453] = 10'b1111110111;
mem2[14454] = 10'b1111110111;
mem2[14455] = 10'b1111110111;
mem2[14456] = 10'b1111110111;
mem2[14457] = 10'b1111110111;
mem2[14458] = 10'b1111110111;
mem2[14459] = 10'b1111110111;
mem2[14460] = 10'b1111110111;
mem2[14461] = 10'b1111110111;
mem2[14462] = 10'b1111110111;
mem2[14463] = 10'b1111110111;
mem2[14464] = 10'b1111110111;
mem2[14465] = 10'b1111110111;
mem2[14466] = 10'b1111110111;
mem2[14467] = 10'b1111110111;
mem2[14468] = 10'b1111110111;
mem2[14469] = 10'b1111110111;
mem2[14470] = 10'b1111110111;
mem2[14471] = 10'b1111110111;
mem2[14472] = 10'b1111110111;
mem2[14473] = 10'b1111110111;
mem2[14474] = 10'b1111110111;
mem2[14475] = 10'b1111110111;
mem2[14476] = 10'b1111110111;
mem2[14477] = 10'b1111110111;
mem2[14478] = 10'b1111110111;
mem2[14479] = 10'b1111110111;
mem2[14480] = 10'b1111110111;
mem2[14481] = 10'b1111110111;
mem2[14482] = 10'b1111110111;
mem2[14483] = 10'b1111110111;
mem2[14484] = 10'b1111110111;
mem2[14485] = 10'b1111110111;
mem2[14486] = 10'b1111110111;
mem2[14487] = 10'b1111110111;
mem2[14488] = 10'b1111110111;
mem2[14489] = 10'b1111110111;
mem2[14490] = 10'b1111110111;
mem2[14491] = 10'b1111110111;
mem2[14492] = 10'b1111110111;
mem2[14493] = 10'b1111110111;
mem2[14494] = 10'b1111111000;
mem2[14495] = 10'b1111111000;
mem2[14496] = 10'b1111111000;
mem2[14497] = 10'b1111111000;
mem2[14498] = 10'b1111111000;
mem2[14499] = 10'b1111111000;
mem2[14500] = 10'b1111111000;
mem2[14501] = 10'b1111111000;
mem2[14502] = 10'b1111111000;
mem2[14503] = 10'b1111111000;
mem2[14504] = 10'b1111111000;
mem2[14505] = 10'b1111111000;
mem2[14506] = 10'b1111111000;
mem2[14507] = 10'b1111111000;
mem2[14508] = 10'b1111111000;
mem2[14509] = 10'b1111111000;
mem2[14510] = 10'b1111111000;
mem2[14511] = 10'b1111111000;
mem2[14512] = 10'b1111111000;
mem2[14513] = 10'b1111111000;
mem2[14514] = 10'b1111111000;
mem2[14515] = 10'b1111111000;
mem2[14516] = 10'b1111111000;
mem2[14517] = 10'b1111111000;
mem2[14518] = 10'b1111111000;
mem2[14519] = 10'b1111111000;
mem2[14520] = 10'b1111111000;
mem2[14521] = 10'b1111111000;
mem2[14522] = 10'b1111111000;
mem2[14523] = 10'b1111111000;
mem2[14524] = 10'b1111111000;
mem2[14525] = 10'b1111111000;
mem2[14526] = 10'b1111111000;
mem2[14527] = 10'b1111111000;
mem2[14528] = 10'b1111111000;
mem2[14529] = 10'b1111111000;
mem2[14530] = 10'b1111111000;
mem2[14531] = 10'b1111111000;
mem2[14532] = 10'b1111111000;
mem2[14533] = 10'b1111111000;
mem2[14534] = 10'b1111111000;
mem2[14535] = 10'b1111111000;
mem2[14536] = 10'b1111111000;
mem2[14537] = 10'b1111111000;
mem2[14538] = 10'b1111111000;
mem2[14539] = 10'b1111111000;
mem2[14540] = 10'b1111111000;
mem2[14541] = 10'b1111111000;
mem2[14542] = 10'b1111111000;
mem2[14543] = 10'b1111111000;
mem2[14544] = 10'b1111111000;
mem2[14545] = 10'b1111111000;
mem2[14546] = 10'b1111111000;
mem2[14547] = 10'b1111111000;
mem2[14548] = 10'b1111111000;
mem2[14549] = 10'b1111111000;
mem2[14550] = 10'b1111111001;
mem2[14551] = 10'b1111111001;
mem2[14552] = 10'b1111111001;
mem2[14553] = 10'b1111111001;
mem2[14554] = 10'b1111111001;
mem2[14555] = 10'b1111111001;
mem2[14556] = 10'b1111111001;
mem2[14557] = 10'b1111111001;
mem2[14558] = 10'b1111111001;
mem2[14559] = 10'b1111111001;
mem2[14560] = 10'b1111111001;
mem2[14561] = 10'b1111111001;
mem2[14562] = 10'b1111111001;
mem2[14563] = 10'b1111111001;
mem2[14564] = 10'b1111111001;
mem2[14565] = 10'b1111111001;
mem2[14566] = 10'b1111111001;
mem2[14567] = 10'b1111111001;
mem2[14568] = 10'b1111111001;
mem2[14569] = 10'b1111111001;
mem2[14570] = 10'b1111111001;
mem2[14571] = 10'b1111111001;
mem2[14572] = 10'b1111111001;
mem2[14573] = 10'b1111111001;
mem2[14574] = 10'b1111111001;
mem2[14575] = 10'b1111111001;
mem2[14576] = 10'b1111111001;
mem2[14577] = 10'b1111111001;
mem2[14578] = 10'b1111111001;
mem2[14579] = 10'b1111111001;
mem2[14580] = 10'b1111111001;
mem2[14581] = 10'b1111111001;
mem2[14582] = 10'b1111111001;
mem2[14583] = 10'b1111111001;
mem2[14584] = 10'b1111111001;
mem2[14585] = 10'b1111111001;
mem2[14586] = 10'b1111111001;
mem2[14587] = 10'b1111111001;
mem2[14588] = 10'b1111111001;
mem2[14589] = 10'b1111111001;
mem2[14590] = 10'b1111111001;
mem2[14591] = 10'b1111111001;
mem2[14592] = 10'b1111111001;
mem2[14593] = 10'b1111111001;
mem2[14594] = 10'b1111111001;
mem2[14595] = 10'b1111111001;
mem2[14596] = 10'b1111111001;
mem2[14597] = 10'b1111111001;
mem2[14598] = 10'b1111111001;
mem2[14599] = 10'b1111111001;
mem2[14600] = 10'b1111111001;
mem2[14601] = 10'b1111111001;
mem2[14602] = 10'b1111111001;
mem2[14603] = 10'b1111111001;
mem2[14604] = 10'b1111111001;
mem2[14605] = 10'b1111111001;
mem2[14606] = 10'b1111111001;
mem2[14607] = 10'b1111111001;
mem2[14608] = 10'b1111111001;
mem2[14609] = 10'b1111111001;
mem2[14610] = 10'b1111111001;
mem2[14611] = 10'b1111111010;
mem2[14612] = 10'b1111111010;
mem2[14613] = 10'b1111111010;
mem2[14614] = 10'b1111111010;
mem2[14615] = 10'b1111111010;
mem2[14616] = 10'b1111111010;
mem2[14617] = 10'b1111111010;
mem2[14618] = 10'b1111111010;
mem2[14619] = 10'b1111111010;
mem2[14620] = 10'b1111111010;
mem2[14621] = 10'b1111111010;
mem2[14622] = 10'b1111111010;
mem2[14623] = 10'b1111111010;
mem2[14624] = 10'b1111111010;
mem2[14625] = 10'b1111111010;
mem2[14626] = 10'b1111111010;
mem2[14627] = 10'b1111111010;
mem2[14628] = 10'b1111111010;
mem2[14629] = 10'b1111111010;
mem2[14630] = 10'b1111111010;
mem2[14631] = 10'b1111111010;
mem2[14632] = 10'b1111111010;
mem2[14633] = 10'b1111111010;
mem2[14634] = 10'b1111111010;
mem2[14635] = 10'b1111111010;
mem2[14636] = 10'b1111111010;
mem2[14637] = 10'b1111111010;
mem2[14638] = 10'b1111111010;
mem2[14639] = 10'b1111111010;
mem2[14640] = 10'b1111111010;
mem2[14641] = 10'b1111111010;
mem2[14642] = 10'b1111111010;
mem2[14643] = 10'b1111111010;
mem2[14644] = 10'b1111111010;
mem2[14645] = 10'b1111111010;
mem2[14646] = 10'b1111111010;
mem2[14647] = 10'b1111111010;
mem2[14648] = 10'b1111111010;
mem2[14649] = 10'b1111111010;
mem2[14650] = 10'b1111111010;
mem2[14651] = 10'b1111111010;
mem2[14652] = 10'b1111111010;
mem2[14653] = 10'b1111111010;
mem2[14654] = 10'b1111111010;
mem2[14655] = 10'b1111111010;
mem2[14656] = 10'b1111111010;
mem2[14657] = 10'b1111111010;
mem2[14658] = 10'b1111111010;
mem2[14659] = 10'b1111111010;
mem2[14660] = 10'b1111111010;
mem2[14661] = 10'b1111111010;
mem2[14662] = 10'b1111111010;
mem2[14663] = 10'b1111111010;
mem2[14664] = 10'b1111111010;
mem2[14665] = 10'b1111111010;
mem2[14666] = 10'b1111111010;
mem2[14667] = 10'b1111111010;
mem2[14668] = 10'b1111111010;
mem2[14669] = 10'b1111111010;
mem2[14670] = 10'b1111111010;
mem2[14671] = 10'b1111111010;
mem2[14672] = 10'b1111111010;
mem2[14673] = 10'b1111111010;
mem2[14674] = 10'b1111111010;
mem2[14675] = 10'b1111111010;
mem2[14676] = 10'b1111111011;
mem2[14677] = 10'b1111111011;
mem2[14678] = 10'b1111111011;
mem2[14679] = 10'b1111111011;
mem2[14680] = 10'b1111111011;
mem2[14681] = 10'b1111111011;
mem2[14682] = 10'b1111111011;
mem2[14683] = 10'b1111111011;
mem2[14684] = 10'b1111111011;
mem2[14685] = 10'b1111111011;
mem2[14686] = 10'b1111111011;
mem2[14687] = 10'b1111111011;
mem2[14688] = 10'b1111111011;
mem2[14689] = 10'b1111111011;
mem2[14690] = 10'b1111111011;
mem2[14691] = 10'b1111111011;
mem2[14692] = 10'b1111111011;
mem2[14693] = 10'b1111111011;
mem2[14694] = 10'b1111111011;
mem2[14695] = 10'b1111111011;
mem2[14696] = 10'b1111111011;
mem2[14697] = 10'b1111111011;
mem2[14698] = 10'b1111111011;
mem2[14699] = 10'b1111111011;
mem2[14700] = 10'b1111111011;
mem2[14701] = 10'b1111111011;
mem2[14702] = 10'b1111111011;
mem2[14703] = 10'b1111111011;
mem2[14704] = 10'b1111111011;
mem2[14705] = 10'b1111111011;
mem2[14706] = 10'b1111111011;
mem2[14707] = 10'b1111111011;
mem2[14708] = 10'b1111111011;
mem2[14709] = 10'b1111111011;
mem2[14710] = 10'b1111111011;
mem2[14711] = 10'b1111111011;
mem2[14712] = 10'b1111111011;
mem2[14713] = 10'b1111111011;
mem2[14714] = 10'b1111111011;
mem2[14715] = 10'b1111111011;
mem2[14716] = 10'b1111111011;
mem2[14717] = 10'b1111111011;
mem2[14718] = 10'b1111111011;
mem2[14719] = 10'b1111111011;
mem2[14720] = 10'b1111111011;
mem2[14721] = 10'b1111111011;
mem2[14722] = 10'b1111111011;
mem2[14723] = 10'b1111111011;
mem2[14724] = 10'b1111111011;
mem2[14725] = 10'b1111111011;
mem2[14726] = 10'b1111111011;
mem2[14727] = 10'b1111111011;
mem2[14728] = 10'b1111111011;
mem2[14729] = 10'b1111111011;
mem2[14730] = 10'b1111111011;
mem2[14731] = 10'b1111111011;
mem2[14732] = 10'b1111111011;
mem2[14733] = 10'b1111111011;
mem2[14734] = 10'b1111111011;
mem2[14735] = 10'b1111111011;
mem2[14736] = 10'b1111111011;
mem2[14737] = 10'b1111111011;
mem2[14738] = 10'b1111111011;
mem2[14739] = 10'b1111111011;
mem2[14740] = 10'b1111111011;
mem2[14741] = 10'b1111111011;
mem2[14742] = 10'b1111111011;
mem2[14743] = 10'b1111111011;
mem2[14744] = 10'b1111111011;
mem2[14745] = 10'b1111111011;
mem2[14746] = 10'b1111111011;
mem2[14747] = 10'b1111111011;
mem2[14748] = 10'b1111111100;
mem2[14749] = 10'b1111111100;
mem2[14750] = 10'b1111111100;
mem2[14751] = 10'b1111111100;
mem2[14752] = 10'b1111111100;
mem2[14753] = 10'b1111111100;
mem2[14754] = 10'b1111111100;
mem2[14755] = 10'b1111111100;
mem2[14756] = 10'b1111111100;
mem2[14757] = 10'b1111111100;
mem2[14758] = 10'b1111111100;
mem2[14759] = 10'b1111111100;
mem2[14760] = 10'b1111111100;
mem2[14761] = 10'b1111111100;
mem2[14762] = 10'b1111111100;
mem2[14763] = 10'b1111111100;
mem2[14764] = 10'b1111111100;
mem2[14765] = 10'b1111111100;
mem2[14766] = 10'b1111111100;
mem2[14767] = 10'b1111111100;
mem2[14768] = 10'b1111111100;
mem2[14769] = 10'b1111111100;
mem2[14770] = 10'b1111111100;
mem2[14771] = 10'b1111111100;
mem2[14772] = 10'b1111111100;
mem2[14773] = 10'b1111111100;
mem2[14774] = 10'b1111111100;
mem2[14775] = 10'b1111111100;
mem2[14776] = 10'b1111111100;
mem2[14777] = 10'b1111111100;
mem2[14778] = 10'b1111111100;
mem2[14779] = 10'b1111111100;
mem2[14780] = 10'b1111111100;
mem2[14781] = 10'b1111111100;
mem2[14782] = 10'b1111111100;
mem2[14783] = 10'b1111111100;
mem2[14784] = 10'b1111111100;
mem2[14785] = 10'b1111111100;
mem2[14786] = 10'b1111111100;
mem2[14787] = 10'b1111111100;
mem2[14788] = 10'b1111111100;
mem2[14789] = 10'b1111111100;
mem2[14790] = 10'b1111111100;
mem2[14791] = 10'b1111111100;
mem2[14792] = 10'b1111111100;
mem2[14793] = 10'b1111111100;
mem2[14794] = 10'b1111111100;
mem2[14795] = 10'b1111111100;
mem2[14796] = 10'b1111111100;
mem2[14797] = 10'b1111111100;
mem2[14798] = 10'b1111111100;
mem2[14799] = 10'b1111111100;
mem2[14800] = 10'b1111111100;
mem2[14801] = 10'b1111111100;
mem2[14802] = 10'b1111111100;
mem2[14803] = 10'b1111111100;
mem2[14804] = 10'b1111111100;
mem2[14805] = 10'b1111111100;
mem2[14806] = 10'b1111111100;
mem2[14807] = 10'b1111111100;
mem2[14808] = 10'b1111111100;
mem2[14809] = 10'b1111111100;
mem2[14810] = 10'b1111111100;
mem2[14811] = 10'b1111111100;
mem2[14812] = 10'b1111111100;
mem2[14813] = 10'b1111111100;
mem2[14814] = 10'b1111111100;
mem2[14815] = 10'b1111111100;
mem2[14816] = 10'b1111111100;
mem2[14817] = 10'b1111111100;
mem2[14818] = 10'b1111111100;
mem2[14819] = 10'b1111111100;
mem2[14820] = 10'b1111111100;
mem2[14821] = 10'b1111111100;
mem2[14822] = 10'b1111111100;
mem2[14823] = 10'b1111111100;
mem2[14824] = 10'b1111111100;
mem2[14825] = 10'b1111111100;
mem2[14826] = 10'b1111111100;
mem2[14827] = 10'b1111111100;
mem2[14828] = 10'b1111111100;
mem2[14829] = 10'b1111111100;
mem2[14830] = 10'b1111111101;
mem2[14831] = 10'b1111111101;
mem2[14832] = 10'b1111111101;
mem2[14833] = 10'b1111111101;
mem2[14834] = 10'b1111111101;
mem2[14835] = 10'b1111111101;
mem2[14836] = 10'b1111111101;
mem2[14837] = 10'b1111111101;
mem2[14838] = 10'b1111111101;
mem2[14839] = 10'b1111111101;
mem2[14840] = 10'b1111111101;
mem2[14841] = 10'b1111111101;
mem2[14842] = 10'b1111111101;
mem2[14843] = 10'b1111111101;
mem2[14844] = 10'b1111111101;
mem2[14845] = 10'b1111111101;
mem2[14846] = 10'b1111111101;
mem2[14847] = 10'b1111111101;
mem2[14848] = 10'b1111111101;
mem2[14849] = 10'b1111111101;
mem2[14850] = 10'b1111111101;
mem2[14851] = 10'b1111111101;
mem2[14852] = 10'b1111111101;
mem2[14853] = 10'b1111111101;
mem2[14854] = 10'b1111111101;
mem2[14855] = 10'b1111111101;
mem2[14856] = 10'b1111111101;
mem2[14857] = 10'b1111111101;
mem2[14858] = 10'b1111111101;
mem2[14859] = 10'b1111111101;
mem2[14860] = 10'b1111111101;
mem2[14861] = 10'b1111111101;
mem2[14862] = 10'b1111111101;
mem2[14863] = 10'b1111111101;
mem2[14864] = 10'b1111111101;
mem2[14865] = 10'b1111111101;
mem2[14866] = 10'b1111111101;
mem2[14867] = 10'b1111111101;
mem2[14868] = 10'b1111111101;
mem2[14869] = 10'b1111111101;
mem2[14870] = 10'b1111111101;
mem2[14871] = 10'b1111111101;
mem2[14872] = 10'b1111111101;
mem2[14873] = 10'b1111111101;
mem2[14874] = 10'b1111111101;
mem2[14875] = 10'b1111111101;
mem2[14876] = 10'b1111111101;
mem2[14877] = 10'b1111111101;
mem2[14878] = 10'b1111111101;
mem2[14879] = 10'b1111111101;
mem2[14880] = 10'b1111111101;
mem2[14881] = 10'b1111111101;
mem2[14882] = 10'b1111111101;
mem2[14883] = 10'b1111111101;
mem2[14884] = 10'b1111111101;
mem2[14885] = 10'b1111111101;
mem2[14886] = 10'b1111111101;
mem2[14887] = 10'b1111111101;
mem2[14888] = 10'b1111111101;
mem2[14889] = 10'b1111111101;
mem2[14890] = 10'b1111111101;
mem2[14891] = 10'b1111111101;
mem2[14892] = 10'b1111111101;
mem2[14893] = 10'b1111111101;
mem2[14894] = 10'b1111111101;
mem2[14895] = 10'b1111111101;
mem2[14896] = 10'b1111111101;
mem2[14897] = 10'b1111111101;
mem2[14898] = 10'b1111111101;
mem2[14899] = 10'b1111111101;
mem2[14900] = 10'b1111111101;
mem2[14901] = 10'b1111111101;
mem2[14902] = 10'b1111111101;
mem2[14903] = 10'b1111111101;
mem2[14904] = 10'b1111111101;
mem2[14905] = 10'b1111111101;
mem2[14906] = 10'b1111111101;
mem2[14907] = 10'b1111111101;
mem2[14908] = 10'b1111111101;
mem2[14909] = 10'b1111111101;
mem2[14910] = 10'b1111111101;
mem2[14911] = 10'b1111111101;
mem2[14912] = 10'b1111111101;
mem2[14913] = 10'b1111111101;
mem2[14914] = 10'b1111111101;
mem2[14915] = 10'b1111111101;
mem2[14916] = 10'b1111111101;
mem2[14917] = 10'b1111111101;
mem2[14918] = 10'b1111111101;
mem2[14919] = 10'b1111111101;
mem2[14920] = 10'b1111111101;
mem2[14921] = 10'b1111111101;
mem2[14922] = 10'b1111111101;
mem2[14923] = 10'b1111111101;
mem2[14924] = 10'b1111111101;
mem2[14925] = 10'b1111111101;
mem2[14926] = 10'b1111111101;
mem2[14927] = 10'b1111111110;
mem2[14928] = 10'b1111111110;
mem2[14929] = 10'b1111111110;
mem2[14930] = 10'b1111111110;
mem2[14931] = 10'b1111111110;
mem2[14932] = 10'b1111111110;
mem2[14933] = 10'b1111111110;
mem2[14934] = 10'b1111111110;
mem2[14935] = 10'b1111111110;
mem2[14936] = 10'b1111111110;
mem2[14937] = 10'b1111111110;
mem2[14938] = 10'b1111111110;
mem2[14939] = 10'b1111111110;
mem2[14940] = 10'b1111111110;
mem2[14941] = 10'b1111111110;
mem2[14942] = 10'b1111111110;
mem2[14943] = 10'b1111111110;
mem2[14944] = 10'b1111111110;
mem2[14945] = 10'b1111111110;
mem2[14946] = 10'b1111111110;
mem2[14947] = 10'b1111111110;
mem2[14948] = 10'b1111111110;
mem2[14949] = 10'b1111111110;
mem2[14950] = 10'b1111111110;
mem2[14951] = 10'b1111111110;
mem2[14952] = 10'b1111111110;
mem2[14953] = 10'b1111111110;
mem2[14954] = 10'b1111111110;
mem2[14955] = 10'b1111111110;
mem2[14956] = 10'b1111111110;
mem2[14957] = 10'b1111111110;
mem2[14958] = 10'b1111111110;
mem2[14959] = 10'b1111111110;
mem2[14960] = 10'b1111111110;
mem2[14961] = 10'b1111111110;
mem2[14962] = 10'b1111111110;
mem2[14963] = 10'b1111111110;
mem2[14964] = 10'b1111111110;
mem2[14965] = 10'b1111111110;
mem2[14966] = 10'b1111111110;
mem2[14967] = 10'b1111111110;
mem2[14968] = 10'b1111111110;
mem2[14969] = 10'b1111111110;
mem2[14970] = 10'b1111111110;
mem2[14971] = 10'b1111111110;
mem2[14972] = 10'b1111111110;
mem2[14973] = 10'b1111111110;
mem2[14974] = 10'b1111111110;
mem2[14975] = 10'b1111111110;
mem2[14976] = 10'b1111111110;
mem2[14977] = 10'b1111111110;
mem2[14978] = 10'b1111111110;
mem2[14979] = 10'b1111111110;
mem2[14980] = 10'b1111111110;
mem2[14981] = 10'b1111111110;
mem2[14982] = 10'b1111111110;
mem2[14983] = 10'b1111111110;
mem2[14984] = 10'b1111111110;
mem2[14985] = 10'b1111111110;
mem2[14986] = 10'b1111111110;
mem2[14987] = 10'b1111111110;
mem2[14988] = 10'b1111111110;
mem2[14989] = 10'b1111111110;
mem2[14990] = 10'b1111111110;
mem2[14991] = 10'b1111111110;
mem2[14992] = 10'b1111111110;
mem2[14993] = 10'b1111111110;
mem2[14994] = 10'b1111111110;
mem2[14995] = 10'b1111111110;
mem2[14996] = 10'b1111111110;
mem2[14997] = 10'b1111111110;
mem2[14998] = 10'b1111111110;
mem2[14999] = 10'b1111111110;
mem2[15000] = 10'b1111111110;
mem2[15001] = 10'b1111111110;
mem2[15002] = 10'b1111111110;
mem2[15003] = 10'b1111111110;
mem2[15004] = 10'b1111111110;
mem2[15005] = 10'b1111111110;
mem2[15006] = 10'b1111111110;
mem2[15007] = 10'b1111111110;
mem2[15008] = 10'b1111111110;
mem2[15009] = 10'b1111111110;
mem2[15010] = 10'b1111111110;
mem2[15011] = 10'b1111111110;
mem2[15012] = 10'b1111111110;
mem2[15013] = 10'b1111111110;
mem2[15014] = 10'b1111111110;
mem2[15015] = 10'b1111111110;
mem2[15016] = 10'b1111111110;
mem2[15017] = 10'b1111111110;
mem2[15018] = 10'b1111111110;
mem2[15019] = 10'b1111111110;
mem2[15020] = 10'b1111111110;
mem2[15021] = 10'b1111111110;
mem2[15022] = 10'b1111111110;
mem2[15023] = 10'b1111111110;
mem2[15024] = 10'b1111111110;
mem2[15025] = 10'b1111111110;
mem2[15026] = 10'b1111111110;
mem2[15027] = 10'b1111111110;
mem2[15028] = 10'b1111111110;
mem2[15029] = 10'b1111111110;
mem2[15030] = 10'b1111111110;
mem2[15031] = 10'b1111111110;
mem2[15032] = 10'b1111111110;
mem2[15033] = 10'b1111111110;
mem2[15034] = 10'b1111111110;
mem2[15035] = 10'b1111111110;
mem2[15036] = 10'b1111111110;
mem2[15037] = 10'b1111111110;
mem2[15038] = 10'b1111111110;
mem2[15039] = 10'b1111111110;
mem2[15040] = 10'b1111111110;
mem2[15041] = 10'b1111111110;
mem2[15042] = 10'b1111111110;
mem2[15043] = 10'b1111111110;
mem2[15044] = 10'b1111111110;
mem2[15045] = 10'b1111111110;
mem2[15046] = 10'b1111111110;
mem2[15047] = 10'b1111111110;
mem2[15048] = 10'b1111111110;
mem2[15049] = 10'b1111111110;
mem2[15050] = 10'b1111111110;
mem2[15051] = 10'b1111111110;
mem2[15052] = 10'b1111111110;
mem2[15053] = 10'b1111111110;
mem2[15054] = 10'b1111111111;
mem2[15055] = 10'b1111111111;
mem2[15056] = 10'b1111111111;
mem2[15057] = 10'b1111111111;
mem2[15058] = 10'b1111111111;
mem2[15059] = 10'b1111111111;
mem2[15060] = 10'b1111111111;
mem2[15061] = 10'b1111111111;
mem2[15062] = 10'b1111111111;
mem2[15063] = 10'b1111111111;
mem2[15064] = 10'b1111111111;
mem2[15065] = 10'b1111111111;
mem2[15066] = 10'b1111111111;
mem2[15067] = 10'b1111111111;
mem2[15068] = 10'b1111111111;
mem2[15069] = 10'b1111111111;
mem2[15070] = 10'b1111111111;
mem2[15071] = 10'b1111111111;
mem2[15072] = 10'b1111111111;
mem2[15073] = 10'b1111111111;
mem2[15074] = 10'b1111111111;
mem2[15075] = 10'b1111111111;
mem2[15076] = 10'b1111111111;
mem2[15077] = 10'b1111111111;
mem2[15078] = 10'b1111111111;
mem2[15079] = 10'b1111111111;
mem2[15080] = 10'b1111111111;
mem2[15081] = 10'b1111111111;
mem2[15082] = 10'b1111111111;
mem2[15083] = 10'b1111111111;
mem2[15084] = 10'b1111111111;
mem2[15085] = 10'b1111111111;
mem2[15086] = 10'b1111111111;
mem2[15087] = 10'b1111111111;
mem2[15088] = 10'b1111111111;
mem2[15089] = 10'b1111111111;
mem2[15090] = 10'b1111111111;
mem2[15091] = 10'b1111111111;
mem2[15092] = 10'b1111111111;
mem2[15093] = 10'b1111111111;
mem2[15094] = 10'b1111111111;
mem2[15095] = 10'b1111111111;
mem2[15096] = 10'b1111111111;
mem2[15097] = 10'b1111111111;
mem2[15098] = 10'b1111111111;
mem2[15099] = 10'b1111111111;
mem2[15100] = 10'b1111111111;
mem2[15101] = 10'b1111111111;
mem2[15102] = 10'b1111111111;
mem2[15103] = 10'b1111111111;
mem2[15104] = 10'b1111111111;
mem2[15105] = 10'b1111111111;
mem2[15106] = 10'b1111111111;
mem2[15107] = 10'b1111111111;
mem2[15108] = 10'b1111111111;
mem2[15109] = 10'b1111111111;
mem2[15110] = 10'b1111111111;
mem2[15111] = 10'b1111111111;
mem2[15112] = 10'b1111111111;
mem2[15113] = 10'b1111111111;
mem2[15114] = 10'b1111111111;
mem2[15115] = 10'b1111111111;
mem2[15116] = 10'b1111111111;
mem2[15117] = 10'b1111111111;
mem2[15118] = 10'b1111111111;
mem2[15119] = 10'b1111111111;
mem2[15120] = 10'b1111111111;
mem2[15121] = 10'b1111111111;
mem2[15122] = 10'b1111111111;
mem2[15123] = 10'b1111111111;
mem2[15124] = 10'b1111111111;
mem2[15125] = 10'b1111111111;
mem2[15126] = 10'b1111111111;
mem2[15127] = 10'b1111111111;
mem2[15128] = 10'b1111111111;
mem2[15129] = 10'b1111111111;
mem2[15130] = 10'b1111111111;
mem2[15131] = 10'b1111111111;
mem2[15132] = 10'b1111111111;
mem2[15133] = 10'b1111111111;
mem2[15134] = 10'b1111111111;
mem2[15135] = 10'b1111111111;
mem2[15136] = 10'b1111111111;
mem2[15137] = 10'b1111111111;
mem2[15138] = 10'b1111111111;
mem2[15139] = 10'b1111111111;
mem2[15140] = 10'b1111111111;
mem2[15141] = 10'b1111111111;
mem2[15142] = 10'b1111111111;
mem2[15143] = 10'b1111111111;
mem2[15144] = 10'b1111111111;
mem2[15145] = 10'b1111111111;
mem2[15146] = 10'b1111111111;
mem2[15147] = 10'b1111111111;
mem2[15148] = 10'b1111111111;
mem2[15149] = 10'b1111111111;
mem2[15150] = 10'b1111111111;
mem2[15151] = 10'b1111111111;
mem2[15152] = 10'b1111111111;
mem2[15153] = 10'b1111111111;
mem2[15154] = 10'b1111111111;
mem2[15155] = 10'b1111111111;
mem2[15156] = 10'b1111111111;
mem2[15157] = 10'b1111111111;
mem2[15158] = 10'b1111111111;
mem2[15159] = 10'b1111111111;
mem2[15160] = 10'b1111111111;
mem2[15161] = 10'b1111111111;
mem2[15162] = 10'b1111111111;
mem2[15163] = 10'b1111111111;
mem2[15164] = 10'b1111111111;
mem2[15165] = 10'b1111111111;
mem2[15166] = 10'b1111111111;
mem2[15167] = 10'b1111111111;
mem2[15168] = 10'b1111111111;
mem2[15169] = 10'b1111111111;
mem2[15170] = 10'b1111111111;
mem2[15171] = 10'b1111111111;
mem2[15172] = 10'b1111111111;
mem2[15173] = 10'b1111111111;
mem2[15174] = 10'b1111111111;
mem2[15175] = 10'b1111111111;
mem2[15176] = 10'b1111111111;
mem2[15177] = 10'b1111111111;
mem2[15178] = 10'b1111111111;
mem2[15179] = 10'b1111111111;
mem2[15180] = 10'b1111111111;
mem2[15181] = 10'b1111111111;
mem2[15182] = 10'b1111111111;
mem2[15183] = 10'b1111111111;
mem2[15184] = 10'b1111111111;
mem2[15185] = 10'b1111111111;
mem2[15186] = 10'b1111111111;
mem2[15187] = 10'b1111111111;
mem2[15188] = 10'b1111111111;
mem2[15189] = 10'b1111111111;
mem2[15190] = 10'b1111111111;
mem2[15191] = 10'b1111111111;
mem2[15192] = 10'b1111111111;
mem2[15193] = 10'b1111111111;
mem2[15194] = 10'b1111111111;
mem2[15195] = 10'b1111111111;
mem2[15196] = 10'b1111111111;
mem2[15197] = 10'b1111111111;
mem2[15198] = 10'b1111111111;
mem2[15199] = 10'b1111111111;
mem2[15200] = 10'b1111111111;
mem2[15201] = 10'b1111111111;
mem2[15202] = 10'b1111111111;
mem2[15203] = 10'b1111111111;
mem2[15204] = 10'b1111111111;
mem2[15205] = 10'b1111111111;
mem2[15206] = 10'b1111111111;
mem2[15207] = 10'b1111111111;
mem2[15208] = 10'b1111111111;
mem2[15209] = 10'b1111111111;
mem2[15210] = 10'b1111111111;
mem2[15211] = 10'b1111111111;
mem2[15212] = 10'b1111111111;
mem2[15213] = 10'b1111111111;
mem2[15214] = 10'b1111111111;
mem2[15215] = 10'b1111111111;
mem2[15216] = 10'b1111111111;
mem2[15217] = 10'b1111111111;
mem2[15218] = 10'b1111111111;
mem2[15219] = 10'b1111111111;
mem2[15220] = 10'b1111111111;
mem2[15221] = 10'b1111111111;
mem2[15222] = 10'b1111111111;
mem2[15223] = 10'b1111111111;
mem2[15224] = 10'b1111111111;
mem2[15225] = 10'b1111111111;
mem2[15226] = 10'b1111111111;
mem2[15227] = 10'b1111111111;
mem2[15228] = 10'b1111111111;
mem2[15229] = 10'b1111111111;
mem2[15230] = 10'b1111111111;
mem2[15231] = 10'b1111111111;
mem2[15232] = 10'b1111111111;
mem2[15233] = 10'b1111111111;
mem2[15234] = 10'b1111111111;
mem2[15235] = 10'b1111111111;
mem2[15236] = 10'b1111111111;
mem2[15237] = 10'b1111111111;
mem2[15238] = 10'b1111111111;
mem2[15239] = 10'b1111111111;
mem2[15240] = 10'b1111111111;
mem2[15241] = 10'b1111111111;
mem2[15242] = 10'b1111111111;
mem2[15243] = 10'b1111111111;
mem2[15244] = 10'b1111111111;
mem2[15245] = 10'b1111111111;
mem2[15246] = 10'b1111111111;
mem2[15247] = 10'b1111111111;
mem2[15248] = 10'b1111111111;
mem2[15249] = 10'b1111111111;
mem2[15250] = 10'b1111111111;
mem2[15251] = 10'b1111111111;
mem2[15252] = 10'b1111111111;
mem2[15253] = 10'b1111111111;
mem2[15254] = 10'b1111111111;
mem2[15255] = 10'b1111111111;
mem2[15256] = 10'b1111111111;
mem2[15257] = 10'b1111111111;
mem2[15258] = 10'b1111111111;
mem2[15259] = 10'b1111111111;
mem2[15260] = 10'b1111111111;
mem2[15261] = 10'b1111111111;
mem2[15262] = 10'b1111111111;
mem2[15263] = 10'b1111111111;
mem2[15264] = 10'b1111111111;
mem2[15265] = 10'b1111111111;
mem2[15266] = 10'b1111111111;
mem2[15267] = 10'b1111111111;
mem2[15268] = 10'b1111111111;
mem2[15269] = 10'b1111111111;
mem2[15270] = 10'b1111111111;
mem2[15271] = 10'b1111111111;
mem2[15272] = 10'b1111111111;
mem2[15273] = 10'b1111111111;
mem2[15274] = 10'b1111111111;
mem2[15275] = 10'b1111111111;
mem2[15276] = 10'b1111111111;
mem2[15277] = 10'b1111111111;
mem2[15278] = 10'b1111111111;
mem2[15279] = 10'b1111111111;
mem2[15280] = 10'b1111111111;
mem2[15281] = 10'b1111111111;
mem2[15282] = 10'b1111111111;
mem2[15283] = 10'b1111111111;
mem2[15284] = 10'b1111111111;
mem2[15285] = 10'b1111111111;
mem2[15286] = 10'b1111111111;
mem2[15287] = 10'b1111111111;
mem2[15288] = 10'b1111111111;
mem2[15289] = 10'b1111111111;
mem2[15290] = 10'b1111111111;
mem2[15291] = 10'b1111111111;
mem2[15292] = 10'b1111111111;
mem2[15293] = 10'b1111111111;
mem2[15294] = 10'b1111111111;
mem2[15295] = 10'b1111111111;
mem2[15296] = 10'b1111111111;
mem2[15297] = 10'b1111111111;
mem2[15298] = 10'b1111111111;
mem2[15299] = 10'b1111111111;
mem2[15300] = 10'b1111111111;
mem2[15301] = 10'b1111111111;
mem2[15302] = 10'b1111111111;
mem2[15303] = 10'b1111111111;
mem2[15304] = 10'b1111111111;
mem2[15305] = 10'b1111111111;
mem2[15306] = 10'b1111111111;
mem2[15307] = 10'b1111111111;
mem2[15308] = 10'b1111111111;
mem2[15309] = 10'b1111111111;
mem2[15310] = 10'b1111111111;
mem2[15311] = 10'b1111111111;
mem2[15312] = 10'b1111111111;
mem2[15313] = 10'b1111111111;
mem2[15314] = 10'b1111111111;
mem2[15315] = 10'b1111111111;
mem2[15316] = 10'b1111111111;
mem2[15317] = 10'b1111111111;
mem2[15318] = 10'b1111111111;
mem2[15319] = 10'b1111111111;
mem2[15320] = 10'b1111111111;
mem2[15321] = 10'b1111111111;
mem2[15322] = 10'b1111111111;
mem2[15323] = 10'b1111111111;
mem2[15324] = 10'b1111111111;
mem2[15325] = 10'b1111111111;
mem2[15326] = 10'b1111111111;
mem2[15327] = 10'b1111111111;
mem2[15328] = 10'b1111111111;
mem2[15329] = 10'b1111111111;
mem2[15330] = 10'b1111111111;
mem2[15331] = 10'b1111111111;
mem2[15332] = 10'b1111111111;
mem2[15333] = 10'b1111111111;
mem2[15334] = 10'b1111111111;
mem2[15335] = 10'b1111111111;
mem2[15336] = 10'b1111111111;
mem2[15337] = 10'b1111111111;
mem2[15338] = 10'b1111111111;
mem2[15339] = 10'b1111111111;
mem2[15340] = 10'b1111111111;
mem2[15341] = 10'b1111111111;
mem2[15342] = 10'b1111111111;
mem2[15343] = 10'b1111111111;
mem2[15344] = 10'b1111111111;
mem2[15345] = 10'b1111111111;
mem2[15346] = 10'b1111111111;
mem2[15347] = 10'b1111111111;
mem2[15348] = 10'b1111111111;
mem2[15349] = 10'b1111111111;
mem2[15350] = 10'b1111111111;
mem2[15351] = 10'b1111111111;
mem2[15352] = 10'b1111111111;
mem2[15353] = 10'b1111111111;
mem2[15354] = 10'b1111111111;
mem2[15355] = 10'b1111111111;
mem2[15356] = 10'b1111111111;
mem2[15357] = 10'b1111111111;
mem2[15358] = 10'b1111111111;
mem2[15359] = 10'b1111111111;


end


always @(posedge clk) begin
	output_data_2 =mem2[selector2] ;
end


//assign output_data_2 = mem2[selector2];

endmodule