module mem1(

	input clk1,
	//input reset_mem1,
	input  wire[13:0] selector1,
	output reg[11:0] output_data_1 

);

reg [7:0] mem1 [0:3839];

initial begin
mem1[0] = 8'b00000000;
mem1[1] = 8'b00000000;
mem1[2] = 8'b00000000;
mem1[3] = 8'b00000000;
mem1[4] = 8'b00000000;
mem1[5] = 8'b00000000;
mem1[6] = 8'b00000000;
mem1[7] = 8'b00000000;
mem1[8] = 8'b00000000;
mem1[9] = 8'b00000000;
mem1[10] = 8'b00000000;
mem1[11] = 8'b00000000;
mem1[12] = 8'b00000000;
mem1[13] = 8'b00000000;
mem1[14] = 8'b00000000;
mem1[15] = 8'b00000000;
mem1[16] = 8'b00000000;
mem1[17] = 8'b00000000;
mem1[18] = 8'b00000000;
mem1[19] = 8'b00000000;
mem1[20] = 8'b00000000;
mem1[21] = 8'b00000000;
mem1[22] = 8'b00000000;
mem1[23] = 8'b00000000;
mem1[24] = 8'b00000000;
mem1[25] = 8'b00000000;
mem1[26] = 8'b00000000;
mem1[27] = 8'b00000000;
mem1[28] = 8'b00000000;
mem1[29] = 8'b00000000;
mem1[30] = 8'b00000000;
mem1[31] = 8'b00000000;
mem1[32] = 8'b00000000;
mem1[33] = 8'b00000000;
mem1[34] = 8'b00000000;
mem1[35] = 8'b00000000;
mem1[36] = 8'b00000000;
mem1[37] = 8'b00000000;
mem1[38] = 8'b00000000;
mem1[39] = 8'b00000000;
mem1[40] = 8'b00000000;
mem1[41] = 8'b00000000;
mem1[42] = 8'b00000000;
mem1[43] = 8'b00000000;
mem1[44] = 8'b00000000;
mem1[45] = 8'b00000000;
mem1[46] = 8'b00000000;
mem1[47] = 8'b00000000;
mem1[48] = 8'b00000000;
mem1[49] = 8'b00000000;
mem1[50] = 8'b00000000;
mem1[51] = 8'b00000000;
mem1[52] = 8'b00000000;
mem1[53] = 8'b00000000;
mem1[54] = 8'b00000000;
mem1[55] = 8'b00000000;
mem1[56] = 8'b00000000;
mem1[57] = 8'b00000000;
mem1[58] = 8'b00000000;
mem1[59] = 8'b00000000;
mem1[60] = 8'b00000000;
mem1[61] = 8'b00000000;
mem1[62] = 8'b00000000;
mem1[63] = 8'b00000000;
mem1[64] = 8'b00000000;
mem1[65] = 8'b00000000;
mem1[66] = 8'b00000000;
mem1[67] = 8'b00000000;
mem1[68] = 8'b00000000;
mem1[69] = 8'b00000000;
mem1[70] = 8'b00000000;
mem1[71] = 8'b00000000;
mem1[72] = 8'b00000000;
mem1[73] = 8'b00000000;
mem1[74] = 8'b00000000;
mem1[75] = 8'b00000000;
mem1[76] = 8'b00000000;
mem1[77] = 8'b00000000;
mem1[78] = 8'b00000000;
mem1[79] = 8'b00000000;
mem1[80] = 8'b00000000;
mem1[81] = 8'b00000000;
mem1[82] = 8'b00000000;
mem1[83] = 8'b00000000;
mem1[84] = 8'b00000000;
mem1[85] = 8'b00000000;
mem1[86] = 8'b00000000;
mem1[87] = 8'b00000000;
mem1[88] = 8'b00000000;
mem1[89] = 8'b00000000;
mem1[90] = 8'b00000000;
mem1[91] = 8'b00000000;
mem1[92] = 8'b00000000;
mem1[93] = 8'b00000000;
mem1[94] = 8'b00000000;
mem1[95] = 8'b00000000;
mem1[96] = 8'b00000000;
mem1[97] = 8'b00000000;
mem1[98] = 8'b00000000;
mem1[99] = 8'b00000000;
mem1[100] = 8'b00000000;
mem1[101] = 8'b00000000;
mem1[102] = 8'b00000000;
mem1[103] = 8'b00000000;
mem1[104] = 8'b00000000;
mem1[105] = 8'b00000000;
mem1[106] = 8'b00000000;
mem1[107] = 8'b00000000;
mem1[108] = 8'b00000000;
mem1[109] = 8'b00000000;
mem1[110] = 8'b00000000;
mem1[111] = 8'b00000000;
mem1[112] = 8'b00000000;
mem1[113] = 8'b00000000;
mem1[114] = 8'b00000000;
mem1[115] = 8'b00000000;
mem1[116] = 8'b00000000;
mem1[117] = 8'b00000000;
mem1[118] = 8'b00000000;
mem1[119] = 8'b00000000;
mem1[120] = 8'b00000000;
mem1[121] = 8'b00000000;
mem1[122] = 8'b00000000;
mem1[123] = 8'b00000000;
mem1[124] = 8'b00000000;
mem1[125] = 8'b00000000;
mem1[126] = 8'b00000000;
mem1[127] = 8'b00000000;
mem1[128] = 8'b00000000;
mem1[129] = 8'b00000000;
mem1[130] = 8'b00000000;
mem1[131] = 8'b00000000;
mem1[132] = 8'b00000000;
mem1[133] = 8'b00000000;
mem1[134] = 8'b00000000;
mem1[135] = 8'b00000000;
mem1[136] = 8'b00000000;
mem1[137] = 8'b00000000;
mem1[138] = 8'b00000000;
mem1[139] = 8'b00000000;
mem1[140] = 8'b00000000;
mem1[141] = 8'b00000000;
mem1[142] = 8'b00000000;
mem1[143] = 8'b00000000;
mem1[144] = 8'b00000000;
mem1[145] = 8'b00000000;
mem1[146] = 8'b00000000;
mem1[147] = 8'b00000000;
mem1[148] = 8'b00000000;
mem1[149] = 8'b00000000;
mem1[150] = 8'b00000000;
mem1[151] = 8'b00000000;
mem1[152] = 8'b00000000;
mem1[153] = 8'b00000001;
mem1[154] = 8'b00000001;
mem1[155] = 8'b00000001;
mem1[156] = 8'b00000001;
mem1[157] = 8'b00000001;
mem1[158] = 8'b00000001;
mem1[159] = 8'b00000001;
mem1[160] = 8'b00000001;
mem1[161] = 8'b00000001;
mem1[162] = 8'b00000001;
mem1[163] = 8'b00000001;
mem1[164] = 8'b00000001;
mem1[165] = 8'b00000001;
mem1[166] = 8'b00000001;
mem1[167] = 8'b00000001;
mem1[168] = 8'b00000001;
mem1[169] = 8'b00000001;
mem1[170] = 8'b00000001;
mem1[171] = 8'b00000001;
mem1[172] = 8'b00000001;
mem1[173] = 8'b00000001;
mem1[174] = 8'b00000001;
mem1[175] = 8'b00000001;
mem1[176] = 8'b00000001;
mem1[177] = 8'b00000001;
mem1[178] = 8'b00000001;
mem1[179] = 8'b00000001;
mem1[180] = 8'b00000001;
mem1[181] = 8'b00000001;
mem1[182] = 8'b00000001;
mem1[183] = 8'b00000001;
mem1[184] = 8'b00000001;
mem1[185] = 8'b00000001;
mem1[186] = 8'b00000001;
mem1[187] = 8'b00000001;
mem1[188] = 8'b00000001;
mem1[189] = 8'b00000001;
mem1[190] = 8'b00000001;
mem1[191] = 8'b00000001;
mem1[192] = 8'b00000001;
mem1[193] = 8'b00000001;
mem1[194] = 8'b00000001;
mem1[195] = 8'b00000001;
mem1[196] = 8'b00000001;
mem1[197] = 8'b00000001;
mem1[198] = 8'b00000001;
mem1[199] = 8'b00000001;
mem1[200] = 8'b00000001;
mem1[201] = 8'b00000001;
mem1[202] = 8'b00000001;
mem1[203] = 8'b00000001;
mem1[204] = 8'b00000001;
mem1[205] = 8'b00000001;
mem1[206] = 8'b00000001;
mem1[207] = 8'b00000001;
mem1[208] = 8'b00000001;
mem1[209] = 8'b00000001;
mem1[210] = 8'b00000001;
mem1[211] = 8'b00000001;
mem1[212] = 8'b00000001;
mem1[213] = 8'b00000001;
mem1[214] = 8'b00000001;
mem1[215] = 8'b00000001;
mem1[216] = 8'b00000001;
mem1[217] = 8'b00000010;
mem1[218] = 8'b00000010;
mem1[219] = 8'b00000010;
mem1[220] = 8'b00000010;
mem1[221] = 8'b00000010;
mem1[222] = 8'b00000010;
mem1[223] = 8'b00000010;
mem1[224] = 8'b00000010;
mem1[225] = 8'b00000010;
mem1[226] = 8'b00000010;
mem1[227] = 8'b00000010;
mem1[228] = 8'b00000010;
mem1[229] = 8'b00000010;
mem1[230] = 8'b00000010;
mem1[231] = 8'b00000010;
mem1[232] = 8'b00000010;
mem1[233] = 8'b00000010;
mem1[234] = 8'b00000010;
mem1[235] = 8'b00000010;
mem1[236] = 8'b00000010;
mem1[237] = 8'b00000010;
mem1[238] = 8'b00000010;
mem1[239] = 8'b00000010;
mem1[240] = 8'b00000010;
mem1[241] = 8'b00000010;
mem1[242] = 8'b00000010;
mem1[243] = 8'b00000010;
mem1[244] = 8'b00000010;
mem1[245] = 8'b00000010;
mem1[246] = 8'b00000010;
mem1[247] = 8'b00000010;
mem1[248] = 8'b00000010;
mem1[249] = 8'b00000010;
mem1[250] = 8'b00000010;
mem1[251] = 8'b00000010;
mem1[252] = 8'b00000010;
mem1[253] = 8'b00000010;
mem1[254] = 8'b00000010;
mem1[255] = 8'b00000010;
mem1[256] = 8'b00000010;
mem1[257] = 8'b00000010;
mem1[258] = 8'b00000010;
mem1[259] = 8'b00000010;
mem1[260] = 8'b00000010;
mem1[261] = 8'b00000010;
mem1[262] = 8'b00000010;
mem1[263] = 8'b00000010;
mem1[264] = 8'b00000010;
mem1[265] = 8'b00000011;
mem1[266] = 8'b00000011;
mem1[267] = 8'b00000011;
mem1[268] = 8'b00000011;
mem1[269] = 8'b00000011;
mem1[270] = 8'b00000011;
mem1[271] = 8'b00000011;
mem1[272] = 8'b00000011;
mem1[273] = 8'b00000011;
mem1[274] = 8'b00000011;
mem1[275] = 8'b00000011;
mem1[276] = 8'b00000011;
mem1[277] = 8'b00000011;
mem1[278] = 8'b00000011;
mem1[279] = 8'b00000011;
mem1[280] = 8'b00000011;
mem1[281] = 8'b00000011;
mem1[282] = 8'b00000011;
mem1[283] = 8'b00000011;
mem1[284] = 8'b00000011;
mem1[285] = 8'b00000011;
mem1[286] = 8'b00000011;
mem1[287] = 8'b00000011;
mem1[288] = 8'b00000011;
mem1[289] = 8'b00000011;
mem1[290] = 8'b00000011;
mem1[291] = 8'b00000011;
mem1[292] = 8'b00000011;
mem1[293] = 8'b00000011;
mem1[294] = 8'b00000011;
mem1[295] = 8'b00000011;
mem1[296] = 8'b00000011;
mem1[297] = 8'b00000011;
mem1[298] = 8'b00000011;
mem1[299] = 8'b00000011;
mem1[300] = 8'b00000011;
mem1[301] = 8'b00000011;
mem1[302] = 8'b00000011;
mem1[303] = 8'b00000011;
mem1[304] = 8'b00000011;
mem1[305] = 8'b00000011;
mem1[306] = 8'b00000011;
mem1[307] = 8'b00000100;
mem1[308] = 8'b00000100;
mem1[309] = 8'b00000100;
mem1[310] = 8'b00000100;
mem1[311] = 8'b00000100;
mem1[312] = 8'b00000100;
mem1[313] = 8'b00000100;
mem1[314] = 8'b00000100;
mem1[315] = 8'b00000100;
mem1[316] = 8'b00000100;
mem1[317] = 8'b00000100;
mem1[318] = 8'b00000100;
mem1[319] = 8'b00000100;
mem1[320] = 8'b00000100;
mem1[321] = 8'b00000100;
mem1[322] = 8'b00000100;
mem1[323] = 8'b00000100;
mem1[324] = 8'b00000100;
mem1[325] = 8'b00000100;
mem1[326] = 8'b00000100;
mem1[327] = 8'b00000100;
mem1[328] = 8'b00000100;
mem1[329] = 8'b00000100;
mem1[330] = 8'b00000100;
mem1[331] = 8'b00000100;
mem1[332] = 8'b00000100;
mem1[333] = 8'b00000100;
mem1[334] = 8'b00000100;
mem1[335] = 8'b00000100;
mem1[336] = 8'b00000100;
mem1[337] = 8'b00000100;
mem1[338] = 8'b00000100;
mem1[339] = 8'b00000100;
mem1[340] = 8'b00000100;
mem1[341] = 8'b00000100;
mem1[342] = 8'b00000100;
mem1[343] = 8'b00000101;
mem1[344] = 8'b00000101;
mem1[345] = 8'b00000101;
mem1[346] = 8'b00000101;
mem1[347] = 8'b00000101;
mem1[348] = 8'b00000101;
mem1[349] = 8'b00000101;
mem1[350] = 8'b00000101;
mem1[351] = 8'b00000101;
mem1[352] = 8'b00000101;
mem1[353] = 8'b00000101;
mem1[354] = 8'b00000101;
mem1[355] = 8'b00000101;
mem1[356] = 8'b00000101;
mem1[357] = 8'b00000101;
mem1[358] = 8'b00000101;
mem1[359] = 8'b00000101;
mem1[360] = 8'b00000101;
mem1[361] = 8'b00000101;
mem1[362] = 8'b00000101;
mem1[363] = 8'b00000101;
mem1[364] = 8'b00000101;
mem1[365] = 8'b00000101;
mem1[366] = 8'b00000101;
mem1[367] = 8'b00000101;
mem1[368] = 8'b00000101;
mem1[369] = 8'b00000101;
mem1[370] = 8'b00000101;
mem1[371] = 8'b00000101;
mem1[372] = 8'b00000101;
mem1[373] = 8'b00000101;
mem1[374] = 8'b00000101;
mem1[375] = 8'b00000101;
mem1[376] = 8'b00000110;
mem1[377] = 8'b00000110;
mem1[378] = 8'b00000110;
mem1[379] = 8'b00000110;
mem1[380] = 8'b00000110;
mem1[381] = 8'b00000110;
mem1[382] = 8'b00000110;
mem1[383] = 8'b00000110;
mem1[384] = 8'b00000110;
mem1[385] = 8'b00000110;
mem1[386] = 8'b00000110;
mem1[387] = 8'b00000110;
mem1[388] = 8'b00000110;
mem1[389] = 8'b00000110;
mem1[390] = 8'b00000110;
mem1[391] = 8'b00000110;
mem1[392] = 8'b00000110;
mem1[393] = 8'b00000110;
mem1[394] = 8'b00000110;
mem1[395] = 8'b00000110;
mem1[396] = 8'b00000110;
mem1[397] = 8'b00000110;
mem1[398] = 8'b00000110;
mem1[399] = 8'b00000110;
mem1[400] = 8'b00000110;
mem1[401] = 8'b00000110;
mem1[402] = 8'b00000110;
mem1[403] = 8'b00000110;
mem1[404] = 8'b00000110;
mem1[405] = 8'b00000110;
mem1[406] = 8'b00000111;
mem1[407] = 8'b00000111;
mem1[408] = 8'b00000111;
mem1[409] = 8'b00000111;
mem1[410] = 8'b00000111;
mem1[411] = 8'b00000111;
mem1[412] = 8'b00000111;
mem1[413] = 8'b00000111;
mem1[414] = 8'b00000111;
mem1[415] = 8'b00000111;
mem1[416] = 8'b00000111;
mem1[417] = 8'b00000111;
mem1[418] = 8'b00000111;
mem1[419] = 8'b00000111;
mem1[420] = 8'b00000111;
mem1[421] = 8'b00000111;
mem1[422] = 8'b00000111;
mem1[423] = 8'b00000111;
mem1[424] = 8'b00000111;
mem1[425] = 8'b00000111;
mem1[426] = 8'b00000111;
mem1[427] = 8'b00000111;
mem1[428] = 8'b00000111;
mem1[429] = 8'b00000111;
mem1[430] = 8'b00000111;
mem1[431] = 8'b00000111;
mem1[432] = 8'b00000111;
mem1[433] = 8'b00000111;
mem1[434] = 8'b00000111;
mem1[435] = 8'b00001000;
mem1[436] = 8'b00001000;
mem1[437] = 8'b00001000;
mem1[438] = 8'b00001000;
mem1[439] = 8'b00001000;
mem1[440] = 8'b00001000;
mem1[441] = 8'b00001000;
mem1[442] = 8'b00001000;
mem1[443] = 8'b00001000;
mem1[444] = 8'b00001000;
mem1[445] = 8'b00001000;
mem1[446] = 8'b00001000;
mem1[447] = 8'b00001000;
mem1[448] = 8'b00001000;
mem1[449] = 8'b00001000;
mem1[450] = 8'b00001000;
mem1[451] = 8'b00001000;
mem1[452] = 8'b00001000;
mem1[453] = 8'b00001000;
mem1[454] = 8'b00001000;
mem1[455] = 8'b00001000;
mem1[456] = 8'b00001000;
mem1[457] = 8'b00001000;
mem1[458] = 8'b00001000;
mem1[459] = 8'b00001000;
mem1[460] = 8'b00001000;
mem1[461] = 8'b00001001;
mem1[462] = 8'b00001001;
mem1[463] = 8'b00001001;
mem1[464] = 8'b00001001;
mem1[465] = 8'b00001001;
mem1[466] = 8'b00001001;
mem1[467] = 8'b00001001;
mem1[468] = 8'b00001001;
mem1[469] = 8'b00001001;
mem1[470] = 8'b00001001;
mem1[471] = 8'b00001001;
mem1[472] = 8'b00001001;
mem1[473] = 8'b00001001;
mem1[474] = 8'b00001001;
mem1[475] = 8'b00001001;
mem1[476] = 8'b00001001;
mem1[477] = 8'b00001001;
mem1[478] = 8'b00001001;
mem1[479] = 8'b00001001;
mem1[480] = 8'b00001001;
mem1[481] = 8'b00001001;
mem1[482] = 8'b00001001;
mem1[483] = 8'b00001001;
mem1[484] = 8'b00001001;
mem1[485] = 8'b00001001;
mem1[486] = 8'b00001001;
mem1[487] = 8'b00001010;
mem1[488] = 8'b00001010;
mem1[489] = 8'b00001010;
mem1[490] = 8'b00001010;
mem1[491] = 8'b00001010;
mem1[492] = 8'b00001010;
mem1[493] = 8'b00001010;
mem1[494] = 8'b00001010;
mem1[495] = 8'b00001010;
mem1[496] = 8'b00001010;
mem1[497] = 8'b00001010;
mem1[498] = 8'b00001010;
mem1[499] = 8'b00001010;
mem1[500] = 8'b00001010;
mem1[501] = 8'b00001010;
mem1[502] = 8'b00001010;
mem1[503] = 8'b00001010;
mem1[504] = 8'b00001010;
mem1[505] = 8'b00001010;
mem1[506] = 8'b00001010;
mem1[507] = 8'b00001010;
mem1[508] = 8'b00001010;
mem1[509] = 8'b00001010;
mem1[510] = 8'b00001010;
mem1[511] = 8'b00001011;
mem1[512] = 8'b00001011;
mem1[513] = 8'b00001011;
mem1[514] = 8'b00001011;
mem1[515] = 8'b00001011;
mem1[516] = 8'b00001011;
mem1[517] = 8'b00001011;
mem1[518] = 8'b00001011;
mem1[519] = 8'b00001011;
mem1[520] = 8'b00001011;
mem1[521] = 8'b00001011;
mem1[522] = 8'b00001011;
mem1[523] = 8'b00001011;
mem1[524] = 8'b00001011;
mem1[525] = 8'b00001011;
mem1[526] = 8'b00001011;
mem1[527] = 8'b00001011;
mem1[528] = 8'b00001011;
mem1[529] = 8'b00001011;
mem1[530] = 8'b00001011;
mem1[531] = 8'b00001011;
mem1[532] = 8'b00001011;
mem1[533] = 8'b00001011;
mem1[534] = 8'b00001100;
mem1[535] = 8'b00001100;
mem1[536] = 8'b00001100;
mem1[537] = 8'b00001100;
mem1[538] = 8'b00001100;
mem1[539] = 8'b00001100;
mem1[540] = 8'b00001100;
mem1[541] = 8'b00001100;
mem1[542] = 8'b00001100;
mem1[543] = 8'b00001100;
mem1[544] = 8'b00001100;
mem1[545] = 8'b00001100;
mem1[546] = 8'b00001100;
mem1[547] = 8'b00001100;
mem1[548] = 8'b00001100;
mem1[549] = 8'b00001100;
mem1[550] = 8'b00001100;
mem1[551] = 8'b00001100;
mem1[552] = 8'b00001100;
mem1[553] = 8'b00001100;
mem1[554] = 8'b00001100;
mem1[555] = 8'b00001100;
mem1[556] = 8'b00001101;
mem1[557] = 8'b00001101;
mem1[558] = 8'b00001101;
mem1[559] = 8'b00001101;
mem1[560] = 8'b00001101;
mem1[561] = 8'b00001101;
mem1[562] = 8'b00001101;
mem1[563] = 8'b00001101;
mem1[564] = 8'b00001101;
mem1[565] = 8'b00001101;
mem1[566] = 8'b00001101;
mem1[567] = 8'b00001101;
mem1[568] = 8'b00001101;
mem1[569] = 8'b00001101;
mem1[570] = 8'b00001101;
mem1[571] = 8'b00001101;
mem1[572] = 8'b00001101;
mem1[573] = 8'b00001101;
mem1[574] = 8'b00001101;
mem1[575] = 8'b00001101;
mem1[576] = 8'b00001101;
mem1[577] = 8'b00001110;
mem1[578] = 8'b00001110;
mem1[579] = 8'b00001110;
mem1[580] = 8'b00001110;
mem1[581] = 8'b00001110;
mem1[582] = 8'b00001110;
mem1[583] = 8'b00001110;
mem1[584] = 8'b00001110;
mem1[585] = 8'b00001110;
mem1[586] = 8'b00001110;
mem1[587] = 8'b00001110;
mem1[588] = 8'b00001110;
mem1[589] = 8'b00001110;
mem1[590] = 8'b00001110;
mem1[591] = 8'b00001110;
mem1[592] = 8'b00001110;
mem1[593] = 8'b00001110;
mem1[594] = 8'b00001110;
mem1[595] = 8'b00001110;
mem1[596] = 8'b00001110;
mem1[597] = 8'b00001110;
mem1[598] = 8'b00001111;
mem1[599] = 8'b00001111;
mem1[600] = 8'b00001111;
mem1[601] = 8'b00001111;
mem1[602] = 8'b00001111;
mem1[603] = 8'b00001111;
mem1[604] = 8'b00001111;
mem1[605] = 8'b00001111;
mem1[606] = 8'b00001111;
mem1[607] = 8'b00001111;
mem1[608] = 8'b00001111;
mem1[609] = 8'b00001111;
mem1[610] = 8'b00001111;
mem1[611] = 8'b00001111;
mem1[612] = 8'b00001111;
mem1[613] = 8'b00001111;
mem1[614] = 8'b00001111;
mem1[615] = 8'b00001111;
mem1[616] = 8'b00001111;
mem1[617] = 8'b00001111;
mem1[618] = 8'b00010000;
mem1[619] = 8'b00010000;
mem1[620] = 8'b00010000;
mem1[621] = 8'b00010000;
mem1[622] = 8'b00010000;
mem1[623] = 8'b00010000;
mem1[624] = 8'b00010000;
mem1[625] = 8'b00010000;
mem1[626] = 8'b00010000;
mem1[627] = 8'b00010000;
mem1[628] = 8'b00010000;
mem1[629] = 8'b00010000;
mem1[630] = 8'b00010000;
mem1[631] = 8'b00010000;
mem1[632] = 8'b00010000;
mem1[633] = 8'b00010000;
mem1[634] = 8'b00010000;
mem1[635] = 8'b00010000;
mem1[636] = 8'b00010000;
mem1[637] = 8'b00010001;
mem1[638] = 8'b00010001;
mem1[639] = 8'b00010001;
mem1[640] = 8'b00010001;
mem1[641] = 8'b00010001;
mem1[642] = 8'b00010001;
mem1[643] = 8'b00010001;
mem1[644] = 8'b00010001;
mem1[645] = 8'b00010001;
mem1[646] = 8'b00010001;
mem1[647] = 8'b00010001;
mem1[648] = 8'b00010001;
mem1[649] = 8'b00010001;
mem1[650] = 8'b00010001;
mem1[651] = 8'b00010001;
mem1[652] = 8'b00010001;
mem1[653] = 8'b00010001;
mem1[654] = 8'b00010001;
mem1[655] = 8'b00010001;
mem1[656] = 8'b00010010;
mem1[657] = 8'b00010010;
mem1[658] = 8'b00010010;
mem1[659] = 8'b00010010;
mem1[660] = 8'b00010010;
mem1[661] = 8'b00010010;
mem1[662] = 8'b00010010;
mem1[663] = 8'b00010010;
mem1[664] = 8'b00010010;
mem1[665] = 8'b00010010;
mem1[666] = 8'b00010010;
mem1[667] = 8'b00010010;
mem1[668] = 8'b00010010;
mem1[669] = 8'b00010010;
mem1[670] = 8'b00010010;
mem1[671] = 8'b00010010;
mem1[672] = 8'b00010010;
mem1[673] = 8'b00010010;
mem1[674] = 8'b00010010;
mem1[675] = 8'b00010011;
mem1[676] = 8'b00010011;
mem1[677] = 8'b00010011;
mem1[678] = 8'b00010011;
mem1[679] = 8'b00010011;
mem1[680] = 8'b00010011;
mem1[681] = 8'b00010011;
mem1[682] = 8'b00010011;
mem1[683] = 8'b00010011;
mem1[684] = 8'b00010011;
mem1[685] = 8'b00010011;
mem1[686] = 8'b00010011;
mem1[687] = 8'b00010011;
mem1[688] = 8'b00010011;
mem1[689] = 8'b00010011;
mem1[690] = 8'b00010011;
mem1[691] = 8'b00010011;
mem1[692] = 8'b00010011;
mem1[693] = 8'b00010100;
mem1[694] = 8'b00010100;
mem1[695] = 8'b00010100;
mem1[696] = 8'b00010100;
mem1[697] = 8'b00010100;
mem1[698] = 8'b00010100;
mem1[699] = 8'b00010100;
mem1[700] = 8'b00010100;
mem1[701] = 8'b00010100;
mem1[702] = 8'b00010100;
mem1[703] = 8'b00010100;
mem1[704] = 8'b00010100;
mem1[705] = 8'b00010100;
mem1[706] = 8'b00010100;
mem1[707] = 8'b00010100;
mem1[708] = 8'b00010100;
mem1[709] = 8'b00010100;
mem1[710] = 8'b00010101;
mem1[711] = 8'b00010101;
mem1[712] = 8'b00010101;
mem1[713] = 8'b00010101;
mem1[714] = 8'b00010101;
mem1[715] = 8'b00010101;
mem1[716] = 8'b00010101;
mem1[717] = 8'b00010101;
mem1[718] = 8'b00010101;
mem1[719] = 8'b00010101;
mem1[720] = 8'b00010101;
mem1[721] = 8'b00010101;
mem1[722] = 8'b00010101;
mem1[723] = 8'b00010101;
mem1[724] = 8'b00010101;
mem1[725] = 8'b00010101;
mem1[726] = 8'b00010101;
mem1[727] = 8'b00010110;
mem1[728] = 8'b00010110;
mem1[729] = 8'b00010110;
mem1[730] = 8'b00010110;
mem1[731] = 8'b00010110;
mem1[732] = 8'b00010110;
mem1[733] = 8'b00010110;
mem1[734] = 8'b00010110;
mem1[735] = 8'b00010110;
mem1[736] = 8'b00010110;
mem1[737] = 8'b00010110;
mem1[738] = 8'b00010110;
mem1[739] = 8'b00010110;
mem1[740] = 8'b00010110;
mem1[741] = 8'b00010110;
mem1[742] = 8'b00010110;
mem1[743] = 8'b00010110;
mem1[744] = 8'b00010111;
mem1[745] = 8'b00010111;
mem1[746] = 8'b00010111;
mem1[747] = 8'b00010111;
mem1[748] = 8'b00010111;
mem1[749] = 8'b00010111;
mem1[750] = 8'b00010111;
mem1[751] = 8'b00010111;
mem1[752] = 8'b00010111;
mem1[753] = 8'b00010111;
mem1[754] = 8'b00010111;
mem1[755] = 8'b00010111;
mem1[756] = 8'b00010111;
mem1[757] = 8'b00010111;
mem1[758] = 8'b00010111;
mem1[759] = 8'b00010111;
mem1[760] = 8'b00010111;
mem1[761] = 8'b00011000;
mem1[762] = 8'b00011000;
mem1[763] = 8'b00011000;
mem1[764] = 8'b00011000;
mem1[765] = 8'b00011000;
mem1[766] = 8'b00011000;
mem1[767] = 8'b00011000;
mem1[768] = 8'b00011000;
mem1[769] = 8'b00011000;
mem1[770] = 8'b00011000;
mem1[771] = 8'b00011000;
mem1[772] = 8'b00011000;
mem1[773] = 8'b00011000;
mem1[774] = 8'b00011000;
mem1[775] = 8'b00011000;
mem1[776] = 8'b00011000;
mem1[777] = 8'b00011001;
mem1[778] = 8'b00011001;
mem1[779] = 8'b00011001;
mem1[780] = 8'b00011001;
mem1[781] = 8'b00011001;
mem1[782] = 8'b00011001;
mem1[783] = 8'b00011001;
mem1[784] = 8'b00011001;
mem1[785] = 8'b00011001;
mem1[786] = 8'b00011001;
mem1[787] = 8'b00011001;
mem1[788] = 8'b00011001;
mem1[789] = 8'b00011001;
mem1[790] = 8'b00011001;
mem1[791] = 8'b00011001;
mem1[792] = 8'b00011001;
mem1[793] = 8'b00011010;
mem1[794] = 8'b00011010;
mem1[795] = 8'b00011010;
mem1[796] = 8'b00011010;
mem1[797] = 8'b00011010;
mem1[798] = 8'b00011010;
mem1[799] = 8'b00011010;
mem1[800] = 8'b00011010;
mem1[801] = 8'b00011010;
mem1[802] = 8'b00011010;
mem1[803] = 8'b00011010;
mem1[804] = 8'b00011010;
mem1[805] = 8'b00011010;
mem1[806] = 8'b00011010;
mem1[807] = 8'b00011010;
mem1[808] = 8'b00011010;
mem1[809] = 8'b00011011;
mem1[810] = 8'b00011011;
mem1[811] = 8'b00011011;
mem1[812] = 8'b00011011;
mem1[813] = 8'b00011011;
mem1[814] = 8'b00011011;
mem1[815] = 8'b00011011;
mem1[816] = 8'b00011011;
mem1[817] = 8'b00011011;
mem1[818] = 8'b00011011;
mem1[819] = 8'b00011011;
mem1[820] = 8'b00011011;
mem1[821] = 8'b00011011;
mem1[822] = 8'b00011011;
mem1[823] = 8'b00011011;
mem1[824] = 8'b00011100;
mem1[825] = 8'b00011100;
mem1[826] = 8'b00011100;
mem1[827] = 8'b00011100;
mem1[828] = 8'b00011100;
mem1[829] = 8'b00011100;
mem1[830] = 8'b00011100;
mem1[831] = 8'b00011100;
mem1[832] = 8'b00011100;
mem1[833] = 8'b00011100;
mem1[834] = 8'b00011100;
mem1[835] = 8'b00011100;
mem1[836] = 8'b00011100;
mem1[837] = 8'b00011100;
mem1[838] = 8'b00011100;
mem1[839] = 8'b00011101;
mem1[840] = 8'b00011101;
mem1[841] = 8'b00011101;
mem1[842] = 8'b00011101;
mem1[843] = 8'b00011101;
mem1[844] = 8'b00011101;
mem1[845] = 8'b00011101;
mem1[846] = 8'b00011101;
mem1[847] = 8'b00011101;
mem1[848] = 8'b00011101;
mem1[849] = 8'b00011101;
mem1[850] = 8'b00011101;
mem1[851] = 8'b00011101;
mem1[852] = 8'b00011101;
mem1[853] = 8'b00011101;
mem1[854] = 8'b00011110;
mem1[855] = 8'b00011110;
mem1[856] = 8'b00011110;
mem1[857] = 8'b00011110;
mem1[858] = 8'b00011110;
mem1[859] = 8'b00011110;
mem1[860] = 8'b00011110;
mem1[861] = 8'b00011110;
mem1[862] = 8'b00011110;
mem1[863] = 8'b00011110;
mem1[864] = 8'b00011110;
mem1[865] = 8'b00011110;
mem1[866] = 8'b00011110;
mem1[867] = 8'b00011110;
mem1[868] = 8'b00011110;
mem1[869] = 8'b00011111;
mem1[870] = 8'b00011111;
mem1[871] = 8'b00011111;
mem1[872] = 8'b00011111;
mem1[873] = 8'b00011111;
mem1[874] = 8'b00011111;
mem1[875] = 8'b00011111;
mem1[876] = 8'b00011111;
mem1[877] = 8'b00011111;
mem1[878] = 8'b00011111;
mem1[879] = 8'b00011111;
mem1[880] = 8'b00011111;
mem1[881] = 8'b00011111;
mem1[882] = 8'b00011111;
mem1[883] = 8'b00011111;
mem1[884] = 8'b00100000;
mem1[885] = 8'b00100000;
mem1[886] = 8'b00100000;
mem1[887] = 8'b00100000;
mem1[888] = 8'b00100000;
mem1[889] = 8'b00100000;
mem1[890] = 8'b00100000;
mem1[891] = 8'b00100000;
mem1[892] = 8'b00100000;
mem1[893] = 8'b00100000;
mem1[894] = 8'b00100000;
mem1[895] = 8'b00100000;
mem1[896] = 8'b00100000;
mem1[897] = 8'b00100000;
mem1[898] = 8'b00100001;
mem1[899] = 8'b00100001;
mem1[900] = 8'b00100001;
mem1[901] = 8'b00100001;
mem1[902] = 8'b00100001;
mem1[903] = 8'b00100001;
mem1[904] = 8'b00100001;
mem1[905] = 8'b00100001;
mem1[906] = 8'b00100001;
mem1[907] = 8'b00100001;
mem1[908] = 8'b00100001;
mem1[909] = 8'b00100001;
mem1[910] = 8'b00100001;
mem1[911] = 8'b00100001;
mem1[912] = 8'b00100010;
mem1[913] = 8'b00100010;
mem1[914] = 8'b00100010;
mem1[915] = 8'b00100010;
mem1[916] = 8'b00100010;
mem1[917] = 8'b00100010;
mem1[918] = 8'b00100010;
mem1[919] = 8'b00100010;
mem1[920] = 8'b00100010;
mem1[921] = 8'b00100010;
mem1[922] = 8'b00100010;
mem1[923] = 8'b00100010;
mem1[924] = 8'b00100010;
mem1[925] = 8'b00100010;
mem1[926] = 8'b00100011;
mem1[927] = 8'b00100011;
mem1[928] = 8'b00100011;
mem1[929] = 8'b00100011;
mem1[930] = 8'b00100011;
mem1[931] = 8'b00100011;
mem1[932] = 8'b00100011;
mem1[933] = 8'b00100011;
mem1[934] = 8'b00100011;
mem1[935] = 8'b00100011;
mem1[936] = 8'b00100011;
mem1[937] = 8'b00100011;
mem1[938] = 8'b00100011;
mem1[939] = 8'b00100011;
mem1[940] = 8'b00100100;
mem1[941] = 8'b00100100;
mem1[942] = 8'b00100100;
mem1[943] = 8'b00100100;
mem1[944] = 8'b00100100;
mem1[945] = 8'b00100100;
mem1[946] = 8'b00100100;
mem1[947] = 8'b00100100;
mem1[948] = 8'b00100100;
mem1[949] = 8'b00100100;
mem1[950] = 8'b00100100;
mem1[951] = 8'b00100100;
mem1[952] = 8'b00100100;
mem1[953] = 8'b00100101;
mem1[954] = 8'b00100101;
mem1[955] = 8'b00100101;
mem1[956] = 8'b00100101;
mem1[957] = 8'b00100101;
mem1[958] = 8'b00100101;
mem1[959] = 8'b00100101;
mem1[960] = 8'b00100101;
mem1[961] = 8'b00100101;
mem1[962] = 8'b00100101;
mem1[963] = 8'b00100101;
mem1[964] = 8'b00100101;
mem1[965] = 8'b00100101;
mem1[966] = 8'b00100101;
mem1[967] = 8'b00100110;
mem1[968] = 8'b00100110;
mem1[969] = 8'b00100110;
mem1[970] = 8'b00100110;
mem1[971] = 8'b00100110;
mem1[972] = 8'b00100110;
mem1[973] = 8'b00100110;
mem1[974] = 8'b00100110;
mem1[975] = 8'b00100110;
mem1[976] = 8'b00100110;
mem1[977] = 8'b00100110;
mem1[978] = 8'b00100110;
mem1[979] = 8'b00100110;
mem1[980] = 8'b00100111;
mem1[981] = 8'b00100111;
mem1[982] = 8'b00100111;
mem1[983] = 8'b00100111;
mem1[984] = 8'b00100111;
mem1[985] = 8'b00100111;
mem1[986] = 8'b00100111;
mem1[987] = 8'b00100111;
mem1[988] = 8'b00100111;
mem1[989] = 8'b00100111;
mem1[990] = 8'b00100111;
mem1[991] = 8'b00100111;
mem1[992] = 8'b00100111;
mem1[993] = 8'b00100111;
mem1[994] = 8'b00101000;
mem1[995] = 8'b00101000;
mem1[996] = 8'b00101000;
mem1[997] = 8'b00101000;
mem1[998] = 8'b00101000;
mem1[999] = 8'b00101000;
mem1[1000] = 8'b00101000;
mem1[1001] = 8'b00101000;
mem1[1002] = 8'b00101000;
mem1[1003] = 8'b00101000;
mem1[1004] = 8'b00101000;
mem1[1005] = 8'b00101000;
mem1[1006] = 8'b00101000;
mem1[1007] = 8'b00101001;
mem1[1008] = 8'b00101001;
mem1[1009] = 8'b00101001;
mem1[1010] = 8'b00101001;
mem1[1011] = 8'b00101001;
mem1[1012] = 8'b00101001;
mem1[1013] = 8'b00101001;
mem1[1014] = 8'b00101001;
mem1[1015] = 8'b00101001;
mem1[1016] = 8'b00101001;
mem1[1017] = 8'b00101001;
mem1[1018] = 8'b00101001;
mem1[1019] = 8'b00101001;
mem1[1020] = 8'b00101010;
mem1[1021] = 8'b00101010;
mem1[1022] = 8'b00101010;
mem1[1023] = 8'b00101010;
mem1[1024] = 8'b00101010;
mem1[1025] = 8'b00101010;
mem1[1026] = 8'b00101010;
mem1[1027] = 8'b00101010;
mem1[1028] = 8'b00101010;
mem1[1029] = 8'b00101010;
mem1[1030] = 8'b00101010;
mem1[1031] = 8'b00101010;
mem1[1032] = 8'b00101011;
mem1[1033] = 8'b00101011;
mem1[1034] = 8'b00101011;
mem1[1035] = 8'b00101011;
mem1[1036] = 8'b00101011;
mem1[1037] = 8'b00101011;
mem1[1038] = 8'b00101011;
mem1[1039] = 8'b00101011;
mem1[1040] = 8'b00101011;
mem1[1041] = 8'b00101011;
mem1[1042] = 8'b00101011;
mem1[1043] = 8'b00101011;
mem1[1044] = 8'b00101011;
mem1[1045] = 8'b00101100;
mem1[1046] = 8'b00101100;
mem1[1047] = 8'b00101100;
mem1[1048] = 8'b00101100;
mem1[1049] = 8'b00101100;
mem1[1050] = 8'b00101100;
mem1[1051] = 8'b00101100;
mem1[1052] = 8'b00101100;
mem1[1053] = 8'b00101100;
mem1[1054] = 8'b00101100;
mem1[1055] = 8'b00101100;
mem1[1056] = 8'b00101100;
mem1[1057] = 8'b00101100;
mem1[1058] = 8'b00101101;
mem1[1059] = 8'b00101101;
mem1[1060] = 8'b00101101;
mem1[1061] = 8'b00101101;
mem1[1062] = 8'b00101101;
mem1[1063] = 8'b00101101;
mem1[1064] = 8'b00101101;
mem1[1065] = 8'b00101101;
mem1[1066] = 8'b00101101;
mem1[1067] = 8'b00101101;
mem1[1068] = 8'b00101101;
mem1[1069] = 8'b00101101;
mem1[1070] = 8'b00101110;
mem1[1071] = 8'b00101110;
mem1[1072] = 8'b00101110;
mem1[1073] = 8'b00101110;
mem1[1074] = 8'b00101110;
mem1[1075] = 8'b00101110;
mem1[1076] = 8'b00101110;
mem1[1077] = 8'b00101110;
mem1[1078] = 8'b00101110;
mem1[1079] = 8'b00101110;
mem1[1080] = 8'b00101110;
mem1[1081] = 8'b00101110;
mem1[1082] = 8'b00101110;
mem1[1083] = 8'b00101111;
mem1[1084] = 8'b00101111;
mem1[1085] = 8'b00101111;
mem1[1086] = 8'b00101111;
mem1[1087] = 8'b00101111;
mem1[1088] = 8'b00101111;
mem1[1089] = 8'b00101111;
mem1[1090] = 8'b00101111;
mem1[1091] = 8'b00101111;
mem1[1092] = 8'b00101111;
mem1[1093] = 8'b00101111;
mem1[1094] = 8'b00101111;
mem1[1095] = 8'b00110000;
mem1[1096] = 8'b00110000;
mem1[1097] = 8'b00110000;
mem1[1098] = 8'b00110000;
mem1[1099] = 8'b00110000;
mem1[1100] = 8'b00110000;
mem1[1101] = 8'b00110000;
mem1[1102] = 8'b00110000;
mem1[1103] = 8'b00110000;
mem1[1104] = 8'b00110000;
mem1[1105] = 8'b00110000;
mem1[1106] = 8'b00110000;
mem1[1107] = 8'b00110001;
mem1[1108] = 8'b00110001;
mem1[1109] = 8'b00110001;
mem1[1110] = 8'b00110001;
mem1[1111] = 8'b00110001;
mem1[1112] = 8'b00110001;
mem1[1113] = 8'b00110001;
mem1[1114] = 8'b00110001;
mem1[1115] = 8'b00110001;
mem1[1116] = 8'b00110001;
mem1[1117] = 8'b00110001;
mem1[1118] = 8'b00110001;
mem1[1119] = 8'b00110010;
mem1[1120] = 8'b00110010;
mem1[1121] = 8'b00110010;
mem1[1122] = 8'b00110010;
mem1[1123] = 8'b00110010;
mem1[1124] = 8'b00110010;
mem1[1125] = 8'b00110010;
mem1[1126] = 8'b00110010;
mem1[1127] = 8'b00110010;
mem1[1128] = 8'b00110010;
mem1[1129] = 8'b00110010;
mem1[1130] = 8'b00110010;
mem1[1131] = 8'b00110011;
mem1[1132] = 8'b00110011;
mem1[1133] = 8'b00110011;
mem1[1134] = 8'b00110011;
mem1[1135] = 8'b00110011;
mem1[1136] = 8'b00110011;
mem1[1137] = 8'b00110011;
mem1[1138] = 8'b00110011;
mem1[1139] = 8'b00110011;
mem1[1140] = 8'b00110011;
mem1[1141] = 8'b00110011;
mem1[1142] = 8'b00110011;
mem1[1143] = 8'b00110100;
mem1[1144] = 8'b00110100;
mem1[1145] = 8'b00110100;
mem1[1146] = 8'b00110100;
mem1[1147] = 8'b00110100;
mem1[1148] = 8'b00110100;
mem1[1149] = 8'b00110100;
mem1[1150] = 8'b00110100;
mem1[1151] = 8'b00110100;
mem1[1152] = 8'b00110100;
mem1[1153] = 8'b00110100;
mem1[1154] = 8'b00110100;
mem1[1155] = 8'b00110101;
mem1[1156] = 8'b00110101;
mem1[1157] = 8'b00110101;
mem1[1158] = 8'b00110101;
mem1[1159] = 8'b00110101;
mem1[1160] = 8'b00110101;
mem1[1161] = 8'b00110101;
mem1[1162] = 8'b00110101;
mem1[1163] = 8'b00110101;
mem1[1164] = 8'b00110101;
mem1[1165] = 8'b00110101;
mem1[1166] = 8'b00110101;
mem1[1167] = 8'b00110110;
mem1[1168] = 8'b00110110;
mem1[1169] = 8'b00110110;
mem1[1170] = 8'b00110110;
mem1[1171] = 8'b00110110;
mem1[1172] = 8'b00110110;
mem1[1173] = 8'b00110110;
mem1[1174] = 8'b00110110;
mem1[1175] = 8'b00110110;
mem1[1176] = 8'b00110110;
mem1[1177] = 8'b00110110;
mem1[1178] = 8'b00110111;
mem1[1179] = 8'b00110111;
mem1[1180] = 8'b00110111;
mem1[1181] = 8'b00110111;
mem1[1182] = 8'b00110111;
mem1[1183] = 8'b00110111;
mem1[1184] = 8'b00110111;
mem1[1185] = 8'b00110111;
mem1[1186] = 8'b00110111;
mem1[1187] = 8'b00110111;
mem1[1188] = 8'b00110111;
mem1[1189] = 8'b00110111;
mem1[1190] = 8'b00111000;
mem1[1191] = 8'b00111000;
mem1[1192] = 8'b00111000;
mem1[1193] = 8'b00111000;
mem1[1194] = 8'b00111000;
mem1[1195] = 8'b00111000;
mem1[1196] = 8'b00111000;
mem1[1197] = 8'b00111000;
mem1[1198] = 8'b00111000;
mem1[1199] = 8'b00111000;
mem1[1200] = 8'b00111000;
mem1[1201] = 8'b00111001;
mem1[1202] = 8'b00111001;
mem1[1203] = 8'b00111001;
mem1[1204] = 8'b00111001;
mem1[1205] = 8'b00111001;
mem1[1206] = 8'b00111001;
mem1[1207] = 8'b00111001;
mem1[1208] = 8'b00111001;
mem1[1209] = 8'b00111001;
mem1[1210] = 8'b00111001;
mem1[1211] = 8'b00111001;
mem1[1212] = 8'b00111001;
mem1[1213] = 8'b00111010;
mem1[1214] = 8'b00111010;
mem1[1215] = 8'b00111010;
mem1[1216] = 8'b00111010;
mem1[1217] = 8'b00111010;
mem1[1218] = 8'b00111010;
mem1[1219] = 8'b00111010;
mem1[1220] = 8'b00111010;
mem1[1221] = 8'b00111010;
mem1[1222] = 8'b00111010;
mem1[1223] = 8'b00111010;
mem1[1224] = 8'b00111011;
mem1[1225] = 8'b00111011;
mem1[1226] = 8'b00111011;
mem1[1227] = 8'b00111011;
mem1[1228] = 8'b00111011;
mem1[1229] = 8'b00111011;
mem1[1230] = 8'b00111011;
mem1[1231] = 8'b00111011;
mem1[1232] = 8'b00111011;
mem1[1233] = 8'b00111011;
mem1[1234] = 8'b00111011;
mem1[1235] = 8'b00111011;
mem1[1236] = 8'b00111100;
mem1[1237] = 8'b00111100;
mem1[1238] = 8'b00111100;
mem1[1239] = 8'b00111100;
mem1[1240] = 8'b00111100;
mem1[1241] = 8'b00111100;
mem1[1242] = 8'b00111100;
mem1[1243] = 8'b00111100;
mem1[1244] = 8'b00111100;
mem1[1245] = 8'b00111100;
mem1[1246] = 8'b00111100;
mem1[1247] = 8'b00111101;
mem1[1248] = 8'b00111101;
mem1[1249] = 8'b00111101;
mem1[1250] = 8'b00111101;
mem1[1251] = 8'b00111101;
mem1[1252] = 8'b00111101;
mem1[1253] = 8'b00111101;
mem1[1254] = 8'b00111101;
mem1[1255] = 8'b00111101;
mem1[1256] = 8'b00111101;
mem1[1257] = 8'b00111101;
mem1[1258] = 8'b00111110;
mem1[1259] = 8'b00111110;
mem1[1260] = 8'b00111110;
mem1[1261] = 8'b00111110;
mem1[1262] = 8'b00111110;
mem1[1263] = 8'b00111110;
mem1[1264] = 8'b00111110;
mem1[1265] = 8'b00111110;
mem1[1266] = 8'b00111110;
mem1[1267] = 8'b00111110;
mem1[1268] = 8'b00111110;
mem1[1269] = 8'b00111111;
mem1[1270] = 8'b00111111;
mem1[1271] = 8'b00111111;
mem1[1272] = 8'b00111111;
mem1[1273] = 8'b00111111;
mem1[1274] = 8'b00111111;
mem1[1275] = 8'b00111111;
mem1[1276] = 8'b00111111;
mem1[1277] = 8'b00111111;
mem1[1278] = 8'b00111111;
mem1[1279] = 8'b00111111;
mem1[1280] = 8'b01000000;
mem1[1281] = 8'b01000000;
mem1[1282] = 8'b01000000;
mem1[1283] = 8'b01000000;
mem1[1284] = 8'b01000000;
mem1[1285] = 8'b01000000;
mem1[1286] = 8'b01000000;
mem1[1287] = 8'b01000000;
mem1[1288] = 8'b01000000;
mem1[1289] = 8'b01000000;
mem1[1290] = 8'b01000000;
mem1[1291] = 8'b01000001;
mem1[1292] = 8'b01000001;
mem1[1293] = 8'b01000001;
mem1[1294] = 8'b01000001;
mem1[1295] = 8'b01000001;
mem1[1296] = 8'b01000001;
mem1[1297] = 8'b01000001;
mem1[1298] = 8'b01000001;
mem1[1299] = 8'b01000001;
mem1[1300] = 8'b01000001;
mem1[1301] = 8'b01000001;
mem1[1302] = 8'b01000010;
mem1[1303] = 8'b01000010;
mem1[1304] = 8'b01000010;
mem1[1305] = 8'b01000010;
mem1[1306] = 8'b01000010;
mem1[1307] = 8'b01000010;
mem1[1308] = 8'b01000010;
mem1[1309] = 8'b01000010;
mem1[1310] = 8'b01000010;
mem1[1311] = 8'b01000010;
mem1[1312] = 8'b01000010;
mem1[1313] = 8'b01000011;
mem1[1314] = 8'b01000011;
mem1[1315] = 8'b01000011;
mem1[1316] = 8'b01000011;
mem1[1317] = 8'b01000011;
mem1[1318] = 8'b01000011;
mem1[1319] = 8'b01000011;
mem1[1320] = 8'b01000011;
mem1[1321] = 8'b01000011;
mem1[1322] = 8'b01000011;
mem1[1323] = 8'b01000011;
mem1[1324] = 8'b01000100;
mem1[1325] = 8'b01000100;
mem1[1326] = 8'b01000100;
mem1[1327] = 8'b01000100;
mem1[1328] = 8'b01000100;
mem1[1329] = 8'b01000100;
mem1[1330] = 8'b01000100;
mem1[1331] = 8'b01000100;
mem1[1332] = 8'b01000100;
mem1[1333] = 8'b01000100;
mem1[1334] = 8'b01000100;
mem1[1335] = 8'b01000101;
mem1[1336] = 8'b01000101;
mem1[1337] = 8'b01000101;
mem1[1338] = 8'b01000101;
mem1[1339] = 8'b01000101;
mem1[1340] = 8'b01000101;
mem1[1341] = 8'b01000101;
mem1[1342] = 8'b01000101;
mem1[1343] = 8'b01000101;
mem1[1344] = 8'b01000101;
mem1[1345] = 8'b01000110;
mem1[1346] = 8'b01000110;
mem1[1347] = 8'b01000110;
mem1[1348] = 8'b01000110;
mem1[1349] = 8'b01000110;
mem1[1350] = 8'b01000110;
mem1[1351] = 8'b01000110;
mem1[1352] = 8'b01000110;
mem1[1353] = 8'b01000110;
mem1[1354] = 8'b01000110;
mem1[1355] = 8'b01000110;
mem1[1356] = 8'b01000111;
mem1[1357] = 8'b01000111;
mem1[1358] = 8'b01000111;
mem1[1359] = 8'b01000111;
mem1[1360] = 8'b01000111;
mem1[1361] = 8'b01000111;
mem1[1362] = 8'b01000111;
mem1[1363] = 8'b01000111;
mem1[1364] = 8'b01000111;
mem1[1365] = 8'b01000111;
mem1[1366] = 8'b01000111;
mem1[1367] = 8'b01001000;
mem1[1368] = 8'b01001000;
mem1[1369] = 8'b01001000;
mem1[1370] = 8'b01001000;
mem1[1371] = 8'b01001000;
mem1[1372] = 8'b01001000;
mem1[1373] = 8'b01001000;
mem1[1374] = 8'b01001000;
mem1[1375] = 8'b01001000;
mem1[1376] = 8'b01001000;
mem1[1377] = 8'b01001001;
mem1[1378] = 8'b01001001;
mem1[1379] = 8'b01001001;
mem1[1380] = 8'b01001001;
mem1[1381] = 8'b01001001;
mem1[1382] = 8'b01001001;
mem1[1383] = 8'b01001001;
mem1[1384] = 8'b01001001;
mem1[1385] = 8'b01001001;
mem1[1386] = 8'b01001001;
mem1[1387] = 8'b01001001;
mem1[1388] = 8'b01001010;
mem1[1389] = 8'b01001010;
mem1[1390] = 8'b01001010;
mem1[1391] = 8'b01001010;
mem1[1392] = 8'b01001010;
mem1[1393] = 8'b01001010;
mem1[1394] = 8'b01001010;
mem1[1395] = 8'b01001010;
mem1[1396] = 8'b01001010;
mem1[1397] = 8'b01001010;
mem1[1398] = 8'b01001011;
mem1[1399] = 8'b01001011;
mem1[1400] = 8'b01001011;
mem1[1401] = 8'b01001011;
mem1[1402] = 8'b01001011;
mem1[1403] = 8'b01001011;
mem1[1404] = 8'b01001011;
mem1[1405] = 8'b01001011;
mem1[1406] = 8'b01001011;
mem1[1407] = 8'b01001011;
mem1[1408] = 8'b01001011;
mem1[1409] = 8'b01001100;
mem1[1410] = 8'b01001100;
mem1[1411] = 8'b01001100;
mem1[1412] = 8'b01001100;
mem1[1413] = 8'b01001100;
mem1[1414] = 8'b01001100;
mem1[1415] = 8'b01001100;
mem1[1416] = 8'b01001100;
mem1[1417] = 8'b01001100;
mem1[1418] = 8'b01001100;
mem1[1419] = 8'b01001101;
mem1[1420] = 8'b01001101;
mem1[1421] = 8'b01001101;
mem1[1422] = 8'b01001101;
mem1[1423] = 8'b01001101;
mem1[1424] = 8'b01001101;
mem1[1425] = 8'b01001101;
mem1[1426] = 8'b01001101;
mem1[1427] = 8'b01001101;
mem1[1428] = 8'b01001101;
mem1[1429] = 8'b01001101;
mem1[1430] = 8'b01001110;
mem1[1431] = 8'b01001110;
mem1[1432] = 8'b01001110;
mem1[1433] = 8'b01001110;
mem1[1434] = 8'b01001110;
mem1[1435] = 8'b01001110;
mem1[1436] = 8'b01001110;
mem1[1437] = 8'b01001110;
mem1[1438] = 8'b01001110;
mem1[1439] = 8'b01001110;
mem1[1440] = 8'b01001111;
mem1[1441] = 8'b01001111;
mem1[1442] = 8'b01001111;
mem1[1443] = 8'b01001111;
mem1[1444] = 8'b01001111;
mem1[1445] = 8'b01001111;
mem1[1446] = 8'b01001111;
mem1[1447] = 8'b01001111;
mem1[1448] = 8'b01001111;
mem1[1449] = 8'b01001111;
mem1[1450] = 8'b01010000;
mem1[1451] = 8'b01010000;
mem1[1452] = 8'b01010000;
mem1[1453] = 8'b01010000;
mem1[1454] = 8'b01010000;
mem1[1455] = 8'b01010000;
mem1[1456] = 8'b01010000;
mem1[1457] = 8'b01010000;
mem1[1458] = 8'b01010000;
mem1[1459] = 8'b01010000;
mem1[1460] = 8'b01010001;
mem1[1461] = 8'b01010001;
mem1[1462] = 8'b01010001;
mem1[1463] = 8'b01010001;
mem1[1464] = 8'b01010001;
mem1[1465] = 8'b01010001;
mem1[1466] = 8'b01010001;
mem1[1467] = 8'b01010001;
mem1[1468] = 8'b01010001;
mem1[1469] = 8'b01010001;
mem1[1470] = 8'b01010001;
mem1[1471] = 8'b01010010;
mem1[1472] = 8'b01010010;
mem1[1473] = 8'b01010010;
mem1[1474] = 8'b01010010;
mem1[1475] = 8'b01010010;
mem1[1476] = 8'b01010010;
mem1[1477] = 8'b01010010;
mem1[1478] = 8'b01010010;
mem1[1479] = 8'b01010010;
mem1[1480] = 8'b01010010;
mem1[1481] = 8'b01010011;
mem1[1482] = 8'b01010011;
mem1[1483] = 8'b01010011;
mem1[1484] = 8'b01010011;
mem1[1485] = 8'b01010011;
mem1[1486] = 8'b01010011;
mem1[1487] = 8'b01010011;
mem1[1488] = 8'b01010011;
mem1[1489] = 8'b01010011;
mem1[1490] = 8'b01010011;
mem1[1491] = 8'b01010100;
mem1[1492] = 8'b01010100;
mem1[1493] = 8'b01010100;
mem1[1494] = 8'b01010100;
mem1[1495] = 8'b01010100;
mem1[1496] = 8'b01010100;
mem1[1497] = 8'b01010100;
mem1[1498] = 8'b01010100;
mem1[1499] = 8'b01010100;
mem1[1500] = 8'b01010100;
mem1[1501] = 8'b01010101;
mem1[1502] = 8'b01010101;
mem1[1503] = 8'b01010101;
mem1[1504] = 8'b01010101;
mem1[1505] = 8'b01010101;
mem1[1506] = 8'b01010101;
mem1[1507] = 8'b01010101;
mem1[1508] = 8'b01010101;
mem1[1509] = 8'b01010101;
mem1[1510] = 8'b01010101;
mem1[1511] = 8'b01010110;
mem1[1512] = 8'b01010110;
mem1[1513] = 8'b01010110;
mem1[1514] = 8'b01010110;
mem1[1515] = 8'b01010110;
mem1[1516] = 8'b01010110;
mem1[1517] = 8'b01010110;
mem1[1518] = 8'b01010110;
mem1[1519] = 8'b01010110;
mem1[1520] = 8'b01010110;
mem1[1521] = 8'b01010110;
mem1[1522] = 8'b01010111;
mem1[1523] = 8'b01010111;
mem1[1524] = 8'b01010111;
mem1[1525] = 8'b01010111;
mem1[1526] = 8'b01010111;
mem1[1527] = 8'b01010111;
mem1[1528] = 8'b01010111;
mem1[1529] = 8'b01010111;
mem1[1530] = 8'b01010111;
mem1[1531] = 8'b01010111;
mem1[1532] = 8'b01011000;
mem1[1533] = 8'b01011000;
mem1[1534] = 8'b01011000;
mem1[1535] = 8'b01011000;
mem1[1536] = 8'b01011000;
mem1[1537] = 8'b01011000;
mem1[1538] = 8'b01011000;
mem1[1539] = 8'b01011000;
mem1[1540] = 8'b01011000;
mem1[1541] = 8'b01011000;
mem1[1542] = 8'b01011001;
mem1[1543] = 8'b01011001;
mem1[1544] = 8'b01011001;
mem1[1545] = 8'b01011001;
mem1[1546] = 8'b01011001;
mem1[1547] = 8'b01011001;
mem1[1548] = 8'b01011001;
mem1[1549] = 8'b01011001;
mem1[1550] = 8'b01011001;
mem1[1551] = 8'b01011001;
mem1[1552] = 8'b01011010;
mem1[1553] = 8'b01011010;
mem1[1554] = 8'b01011010;
mem1[1555] = 8'b01011010;
mem1[1556] = 8'b01011010;
mem1[1557] = 8'b01011010;
mem1[1558] = 8'b01011010;
mem1[1559] = 8'b01011010;
mem1[1560] = 8'b01011010;
mem1[1561] = 8'b01011010;
mem1[1562] = 8'b01011011;
mem1[1563] = 8'b01011011;
mem1[1564] = 8'b01011011;
mem1[1565] = 8'b01011011;
mem1[1566] = 8'b01011011;
mem1[1567] = 8'b01011011;
mem1[1568] = 8'b01011011;
mem1[1569] = 8'b01011011;
mem1[1570] = 8'b01011011;
mem1[1571] = 8'b01011011;
mem1[1572] = 8'b01011100;
mem1[1573] = 8'b01011100;
mem1[1574] = 8'b01011100;
mem1[1575] = 8'b01011100;
mem1[1576] = 8'b01011100;
mem1[1577] = 8'b01011100;
mem1[1578] = 8'b01011100;
mem1[1579] = 8'b01011100;
mem1[1580] = 8'b01011100;
mem1[1581] = 8'b01011100;
mem1[1582] = 8'b01011101;
mem1[1583] = 8'b01011101;
mem1[1584] = 8'b01011101;
mem1[1585] = 8'b01011101;
mem1[1586] = 8'b01011101;
mem1[1587] = 8'b01011101;
mem1[1588] = 8'b01011101;
mem1[1589] = 8'b01011101;
mem1[1590] = 8'b01011101;
mem1[1591] = 8'b01011110;
mem1[1592] = 8'b01011110;
mem1[1593] = 8'b01011110;
mem1[1594] = 8'b01011110;
mem1[1595] = 8'b01011110;
mem1[1596] = 8'b01011110;
mem1[1597] = 8'b01011110;
mem1[1598] = 8'b01011110;
mem1[1599] = 8'b01011110;
mem1[1600] = 8'b01011110;
mem1[1601] = 8'b01011111;
mem1[1602] = 8'b01011111;
mem1[1603] = 8'b01011111;
mem1[1604] = 8'b01011111;
mem1[1605] = 8'b01011111;
mem1[1606] = 8'b01011111;
mem1[1607] = 8'b01011111;
mem1[1608] = 8'b01011111;
mem1[1609] = 8'b01011111;
mem1[1610] = 8'b01011111;
mem1[1611] = 8'b01100000;
mem1[1612] = 8'b01100000;
mem1[1613] = 8'b01100000;
mem1[1614] = 8'b01100000;
mem1[1615] = 8'b01100000;
mem1[1616] = 8'b01100000;
mem1[1617] = 8'b01100000;
mem1[1618] = 8'b01100000;
mem1[1619] = 8'b01100000;
mem1[1620] = 8'b01100000;
mem1[1621] = 8'b01100001;
mem1[1622] = 8'b01100001;
mem1[1623] = 8'b01100001;
mem1[1624] = 8'b01100001;
mem1[1625] = 8'b01100001;
mem1[1626] = 8'b01100001;
mem1[1627] = 8'b01100001;
mem1[1628] = 8'b01100001;
mem1[1629] = 8'b01100001;
mem1[1630] = 8'b01100001;
mem1[1631] = 8'b01100010;
mem1[1632] = 8'b01100010;
mem1[1633] = 8'b01100010;
mem1[1634] = 8'b01100010;
mem1[1635] = 8'b01100010;
mem1[1636] = 8'b01100010;
mem1[1637] = 8'b01100010;
mem1[1638] = 8'b01100010;
mem1[1639] = 8'b01100010;
mem1[1640] = 8'b01100010;
mem1[1641] = 8'b01100011;
mem1[1642] = 8'b01100011;
mem1[1643] = 8'b01100011;
mem1[1644] = 8'b01100011;
mem1[1645] = 8'b01100011;
mem1[1646] = 8'b01100011;
mem1[1647] = 8'b01100011;
mem1[1648] = 8'b01100011;
mem1[1649] = 8'b01100011;
mem1[1650] = 8'b01100100;
mem1[1651] = 8'b01100100;
mem1[1652] = 8'b01100100;
mem1[1653] = 8'b01100100;
mem1[1654] = 8'b01100100;
mem1[1655] = 8'b01100100;
mem1[1656] = 8'b01100100;
mem1[1657] = 8'b01100100;
mem1[1658] = 8'b01100100;
mem1[1659] = 8'b01100100;
mem1[1660] = 8'b01100101;
mem1[1661] = 8'b01100101;
mem1[1662] = 8'b01100101;
mem1[1663] = 8'b01100101;
mem1[1664] = 8'b01100101;
mem1[1665] = 8'b01100101;
mem1[1666] = 8'b01100101;
mem1[1667] = 8'b01100101;
mem1[1668] = 8'b01100101;
mem1[1669] = 8'b01100101;
mem1[1670] = 8'b01100110;
mem1[1671] = 8'b01100110;
mem1[1672] = 8'b01100110;
mem1[1673] = 8'b01100110;
mem1[1674] = 8'b01100110;
mem1[1675] = 8'b01100110;
mem1[1676] = 8'b01100110;
mem1[1677] = 8'b01100110;
mem1[1678] = 8'b01100110;
mem1[1679] = 8'b01100110;
mem1[1680] = 8'b01100111;
mem1[1681] = 8'b01100111;
mem1[1682] = 8'b01100111;
mem1[1683] = 8'b01100111;
mem1[1684] = 8'b01100111;
mem1[1685] = 8'b01100111;
mem1[1686] = 8'b01100111;
mem1[1687] = 8'b01100111;
mem1[1688] = 8'b01100111;
mem1[1689] = 8'b01101000;
mem1[1690] = 8'b01101000;
mem1[1691] = 8'b01101000;
mem1[1692] = 8'b01101000;
mem1[1693] = 8'b01101000;
mem1[1694] = 8'b01101000;
mem1[1695] = 8'b01101000;
mem1[1696] = 8'b01101000;
mem1[1697] = 8'b01101000;
mem1[1698] = 8'b01101000;
mem1[1699] = 8'b01101001;
mem1[1700] = 8'b01101001;
mem1[1701] = 8'b01101001;
mem1[1702] = 8'b01101001;
mem1[1703] = 8'b01101001;
mem1[1704] = 8'b01101001;
mem1[1705] = 8'b01101001;
mem1[1706] = 8'b01101001;
mem1[1707] = 8'b01101001;
mem1[1708] = 8'b01101001;
mem1[1709] = 8'b01101010;
mem1[1710] = 8'b01101010;
mem1[1711] = 8'b01101010;
mem1[1712] = 8'b01101010;
mem1[1713] = 8'b01101010;
mem1[1714] = 8'b01101010;
mem1[1715] = 8'b01101010;
mem1[1716] = 8'b01101010;
mem1[1717] = 8'b01101010;
mem1[1718] = 8'b01101010;
mem1[1719] = 8'b01101011;
mem1[1720] = 8'b01101011;
mem1[1721] = 8'b01101011;
mem1[1722] = 8'b01101011;
mem1[1723] = 8'b01101011;
mem1[1724] = 8'b01101011;
mem1[1725] = 8'b01101011;
mem1[1726] = 8'b01101011;
mem1[1727] = 8'b01101011;
mem1[1728] = 8'b01101100;
mem1[1729] = 8'b01101100;
mem1[1730] = 8'b01101100;
mem1[1731] = 8'b01101100;
mem1[1732] = 8'b01101100;
mem1[1733] = 8'b01101100;
mem1[1734] = 8'b01101100;
mem1[1735] = 8'b01101100;
mem1[1736] = 8'b01101100;
mem1[1737] = 8'b01101100;
mem1[1738] = 8'b01101101;
mem1[1739] = 8'b01101101;
mem1[1740] = 8'b01101101;
mem1[1741] = 8'b01101101;
mem1[1742] = 8'b01101101;
mem1[1743] = 8'b01101101;
mem1[1744] = 8'b01101101;
mem1[1745] = 8'b01101101;
mem1[1746] = 8'b01101101;
mem1[1747] = 8'b01101101;
mem1[1748] = 8'b01101110;
mem1[1749] = 8'b01101110;
mem1[1750] = 8'b01101110;
mem1[1751] = 8'b01101110;
mem1[1752] = 8'b01101110;
mem1[1753] = 8'b01101110;
mem1[1754] = 8'b01101110;
mem1[1755] = 8'b01101110;
mem1[1756] = 8'b01101110;
mem1[1757] = 8'b01101111;
mem1[1758] = 8'b01101111;
mem1[1759] = 8'b01101111;
mem1[1760] = 8'b01101111;
mem1[1761] = 8'b01101111;
mem1[1762] = 8'b01101111;
mem1[1763] = 8'b01101111;
mem1[1764] = 8'b01101111;
mem1[1765] = 8'b01101111;
mem1[1766] = 8'b01101111;
mem1[1767] = 8'b01110000;
mem1[1768] = 8'b01110000;
mem1[1769] = 8'b01110000;
mem1[1770] = 8'b01110000;
mem1[1771] = 8'b01110000;
mem1[1772] = 8'b01110000;
mem1[1773] = 8'b01110000;
mem1[1774] = 8'b01110000;
mem1[1775] = 8'b01110000;
mem1[1776] = 8'b01110001;
mem1[1777] = 8'b01110001;
mem1[1778] = 8'b01110001;
mem1[1779] = 8'b01110001;
mem1[1780] = 8'b01110001;
mem1[1781] = 8'b01110001;
mem1[1782] = 8'b01110001;
mem1[1783] = 8'b01110001;
mem1[1784] = 8'b01110001;
mem1[1785] = 8'b01110001;
mem1[1786] = 8'b01110010;
mem1[1787] = 8'b01110010;
mem1[1788] = 8'b01110010;
mem1[1789] = 8'b01110010;
mem1[1790] = 8'b01110010;
mem1[1791] = 8'b01110010;
mem1[1792] = 8'b01110010;
mem1[1793] = 8'b01110010;
mem1[1794] = 8'b01110010;
mem1[1795] = 8'b01110010;
mem1[1796] = 8'b01110011;
mem1[1797] = 8'b01110011;
mem1[1798] = 8'b01110011;
mem1[1799] = 8'b01110011;
mem1[1800] = 8'b01110011;
mem1[1801] = 8'b01110011;
mem1[1802] = 8'b01110011;
mem1[1803] = 8'b01110011;
mem1[1804] = 8'b01110011;
mem1[1805] = 8'b01110100;
mem1[1806] = 8'b01110100;
mem1[1807] = 8'b01110100;
mem1[1808] = 8'b01110100;
mem1[1809] = 8'b01110100;
mem1[1810] = 8'b01110100;
mem1[1811] = 8'b01110100;
mem1[1812] = 8'b01110100;
mem1[1813] = 8'b01110100;
mem1[1814] = 8'b01110100;
mem1[1815] = 8'b01110101;
mem1[1816] = 8'b01110101;
mem1[1817] = 8'b01110101;
mem1[1818] = 8'b01110101;
mem1[1819] = 8'b01110101;
mem1[1820] = 8'b01110101;
mem1[1821] = 8'b01110101;
mem1[1822] = 8'b01110101;
mem1[1823] = 8'b01110101;
mem1[1824] = 8'b01110110;
mem1[1825] = 8'b01110110;
mem1[1826] = 8'b01110110;
mem1[1827] = 8'b01110110;
mem1[1828] = 8'b01110110;
mem1[1829] = 8'b01110110;
mem1[1830] = 8'b01110110;
mem1[1831] = 8'b01110110;
mem1[1832] = 8'b01110110;
mem1[1833] = 8'b01110110;
mem1[1834] = 8'b01110111;
mem1[1835] = 8'b01110111;
mem1[1836] = 8'b01110111;
mem1[1837] = 8'b01110111;
mem1[1838] = 8'b01110111;
mem1[1839] = 8'b01110111;
mem1[1840] = 8'b01110111;
mem1[1841] = 8'b01110111;
mem1[1842] = 8'b01110111;
mem1[1843] = 8'b01110111;
mem1[1844] = 8'b01111000;
mem1[1845] = 8'b01111000;
mem1[1846] = 8'b01111000;
mem1[1847] = 8'b01111000;
mem1[1848] = 8'b01111000;
mem1[1849] = 8'b01111000;
mem1[1850] = 8'b01111000;
mem1[1851] = 8'b01111000;
mem1[1852] = 8'b01111000;
mem1[1853] = 8'b01111001;
mem1[1854] = 8'b01111001;
mem1[1855] = 8'b01111001;
mem1[1856] = 8'b01111001;
mem1[1857] = 8'b01111001;
mem1[1858] = 8'b01111001;
mem1[1859] = 8'b01111001;
mem1[1860] = 8'b01111001;
mem1[1861] = 8'b01111001;
mem1[1862] = 8'b01111001;
mem1[1863] = 8'b01111010;
mem1[1864] = 8'b01111010;
mem1[1865] = 8'b01111010;
mem1[1866] = 8'b01111010;
mem1[1867] = 8'b01111010;
mem1[1868] = 8'b01111010;
mem1[1869] = 8'b01111010;
mem1[1870] = 8'b01111010;
mem1[1871] = 8'b01111010;
mem1[1872] = 8'b01111011;
mem1[1873] = 8'b01111011;
mem1[1874] = 8'b01111011;
mem1[1875] = 8'b01111011;
mem1[1876] = 8'b01111011;
mem1[1877] = 8'b01111011;
mem1[1878] = 8'b01111011;
mem1[1879] = 8'b01111011;
mem1[1880] = 8'b01111011;
mem1[1881] = 8'b01111011;
mem1[1882] = 8'b01111100;
mem1[1883] = 8'b01111100;
mem1[1884] = 8'b01111100;
mem1[1885] = 8'b01111100;
mem1[1886] = 8'b01111100;
mem1[1887] = 8'b01111100;
mem1[1888] = 8'b01111100;
mem1[1889] = 8'b01111100;
mem1[1890] = 8'b01111100;
mem1[1891] = 8'b01111101;
mem1[1892] = 8'b01111101;
mem1[1893] = 8'b01111101;
mem1[1894] = 8'b01111101;
mem1[1895] = 8'b01111101;
mem1[1896] = 8'b01111101;
mem1[1897] = 8'b01111101;
mem1[1898] = 8'b01111101;
mem1[1899] = 8'b01111101;
mem1[1900] = 8'b01111101;
mem1[1901] = 8'b01111110;
mem1[1902] = 8'b01111110;
mem1[1903] = 8'b01111110;
mem1[1904] = 8'b01111110;
mem1[1905] = 8'b01111110;
mem1[1906] = 8'b01111110;
mem1[1907] = 8'b01111110;
mem1[1908] = 8'b01111110;
mem1[1909] = 8'b01111110;
mem1[1910] = 8'b01111111;
mem1[1911] = 8'b01111111;
mem1[1912] = 8'b01111111;
mem1[1913] = 8'b01111111;
mem1[1914] = 8'b01111111;
mem1[1915] = 8'b01111111;
mem1[1916] = 8'b01111111;
mem1[1917] = 8'b01111111;
mem1[1918] = 8'b01111111;
mem1[1919] = 8'b01111111;
mem1[1920] = 8'b10000000;
mem1[1921] = 8'b10000000;
mem1[1922] = 8'b10000000;
mem1[1923] = 8'b10000000;
mem1[1924] = 8'b10000000;
mem1[1925] = 8'b10000000;
mem1[1926] = 8'b10000000;
mem1[1927] = 8'b10000000;
mem1[1928] = 8'b10000000;
mem1[1929] = 8'b10000000;
mem1[1930] = 8'b10000001;
mem1[1931] = 8'b10000001;
mem1[1932] = 8'b10000001;
mem1[1933] = 8'b10000001;
mem1[1934] = 8'b10000001;
mem1[1935] = 8'b10000001;
mem1[1936] = 8'b10000001;
mem1[1937] = 8'b10000001;
mem1[1938] = 8'b10000001;
mem1[1939] = 8'b10000010;
mem1[1940] = 8'b10000010;
mem1[1941] = 8'b10000010;
mem1[1942] = 8'b10000010;
mem1[1943] = 8'b10000010;
mem1[1944] = 8'b10000010;
mem1[1945] = 8'b10000010;
mem1[1946] = 8'b10000010;
mem1[1947] = 8'b10000010;
mem1[1948] = 8'b10000010;
mem1[1949] = 8'b10000011;
mem1[1950] = 8'b10000011;
mem1[1951] = 8'b10000011;
mem1[1952] = 8'b10000011;
mem1[1953] = 8'b10000011;
mem1[1954] = 8'b10000011;
mem1[1955] = 8'b10000011;
mem1[1956] = 8'b10000011;
mem1[1957] = 8'b10000011;
mem1[1958] = 8'b10000100;
mem1[1959] = 8'b10000100;
mem1[1960] = 8'b10000100;
mem1[1961] = 8'b10000100;
mem1[1962] = 8'b10000100;
mem1[1963] = 8'b10000100;
mem1[1964] = 8'b10000100;
mem1[1965] = 8'b10000100;
mem1[1966] = 8'b10000100;
mem1[1967] = 8'b10000100;
mem1[1968] = 8'b10000101;
mem1[1969] = 8'b10000101;
mem1[1970] = 8'b10000101;
mem1[1971] = 8'b10000101;
mem1[1972] = 8'b10000101;
mem1[1973] = 8'b10000101;
mem1[1974] = 8'b10000101;
mem1[1975] = 8'b10000101;
mem1[1976] = 8'b10000101;
mem1[1977] = 8'b10000110;
mem1[1978] = 8'b10000110;
mem1[1979] = 8'b10000110;
mem1[1980] = 8'b10000110;
mem1[1981] = 8'b10000110;
mem1[1982] = 8'b10000110;
mem1[1983] = 8'b10000110;
mem1[1984] = 8'b10000110;
mem1[1985] = 8'b10000110;
mem1[1986] = 8'b10000110;
mem1[1987] = 8'b10000111;
mem1[1988] = 8'b10000111;
mem1[1989] = 8'b10000111;
mem1[1990] = 8'b10000111;
mem1[1991] = 8'b10000111;
mem1[1992] = 8'b10000111;
mem1[1993] = 8'b10000111;
mem1[1994] = 8'b10000111;
mem1[1995] = 8'b10000111;
mem1[1996] = 8'b10001000;
mem1[1997] = 8'b10001000;
mem1[1998] = 8'b10001000;
mem1[1999] = 8'b10001000;
mem1[2000] = 8'b10001000;
mem1[2001] = 8'b10001000;
mem1[2002] = 8'b10001000;
mem1[2003] = 8'b10001000;
mem1[2004] = 8'b10001000;
mem1[2005] = 8'b10001000;
mem1[2006] = 8'b10001001;
mem1[2007] = 8'b10001001;
mem1[2008] = 8'b10001001;
mem1[2009] = 8'b10001001;
mem1[2010] = 8'b10001001;
mem1[2011] = 8'b10001001;
mem1[2012] = 8'b10001001;
mem1[2013] = 8'b10001001;
mem1[2014] = 8'b10001001;
mem1[2015] = 8'b10001001;
mem1[2016] = 8'b10001010;
mem1[2017] = 8'b10001010;
mem1[2018] = 8'b10001010;
mem1[2019] = 8'b10001010;
mem1[2020] = 8'b10001010;
mem1[2021] = 8'b10001010;
mem1[2022] = 8'b10001010;
mem1[2023] = 8'b10001010;
mem1[2024] = 8'b10001010;
mem1[2025] = 8'b10001011;
mem1[2026] = 8'b10001011;
mem1[2027] = 8'b10001011;
mem1[2028] = 8'b10001011;
mem1[2029] = 8'b10001011;
mem1[2030] = 8'b10001011;
mem1[2031] = 8'b10001011;
mem1[2032] = 8'b10001011;
mem1[2033] = 8'b10001011;
mem1[2034] = 8'b10001011;
mem1[2035] = 8'b10001100;
mem1[2036] = 8'b10001100;
mem1[2037] = 8'b10001100;
mem1[2038] = 8'b10001100;
mem1[2039] = 8'b10001100;
mem1[2040] = 8'b10001100;
mem1[2041] = 8'b10001100;
mem1[2042] = 8'b10001100;
mem1[2043] = 8'b10001100;
mem1[2044] = 8'b10001101;
mem1[2045] = 8'b10001101;
mem1[2046] = 8'b10001101;
mem1[2047] = 8'b10001101;
mem1[2048] = 8'b10001101;
mem1[2049] = 8'b10001101;
mem1[2050] = 8'b10001101;
mem1[2051] = 8'b10001101;
mem1[2052] = 8'b10001101;
mem1[2053] = 8'b10001101;
mem1[2054] = 8'b10001110;
mem1[2055] = 8'b10001110;
mem1[2056] = 8'b10001110;
mem1[2057] = 8'b10001110;
mem1[2058] = 8'b10001110;
mem1[2059] = 8'b10001110;
mem1[2060] = 8'b10001110;
mem1[2061] = 8'b10001110;
mem1[2062] = 8'b10001110;
mem1[2063] = 8'b10001110;
mem1[2064] = 8'b10001111;
mem1[2065] = 8'b10001111;
mem1[2066] = 8'b10001111;
mem1[2067] = 8'b10001111;
mem1[2068] = 8'b10001111;
mem1[2069] = 8'b10001111;
mem1[2070] = 8'b10001111;
mem1[2071] = 8'b10001111;
mem1[2072] = 8'b10001111;
mem1[2073] = 8'b10010000;
mem1[2074] = 8'b10010000;
mem1[2075] = 8'b10010000;
mem1[2076] = 8'b10010000;
mem1[2077] = 8'b10010000;
mem1[2078] = 8'b10010000;
mem1[2079] = 8'b10010000;
mem1[2080] = 8'b10010000;
mem1[2081] = 8'b10010000;
mem1[2082] = 8'b10010000;
mem1[2083] = 8'b10010001;
mem1[2084] = 8'b10010001;
mem1[2085] = 8'b10010001;
mem1[2086] = 8'b10010001;
mem1[2087] = 8'b10010001;
mem1[2088] = 8'b10010001;
mem1[2089] = 8'b10010001;
mem1[2090] = 8'b10010001;
mem1[2091] = 8'b10010001;
mem1[2092] = 8'b10010010;
mem1[2093] = 8'b10010010;
mem1[2094] = 8'b10010010;
mem1[2095] = 8'b10010010;
mem1[2096] = 8'b10010010;
mem1[2097] = 8'b10010010;
mem1[2098] = 8'b10010010;
mem1[2099] = 8'b10010010;
mem1[2100] = 8'b10010010;
mem1[2101] = 8'b10010010;
mem1[2102] = 8'b10010011;
mem1[2103] = 8'b10010011;
mem1[2104] = 8'b10010011;
mem1[2105] = 8'b10010011;
mem1[2106] = 8'b10010011;
mem1[2107] = 8'b10010011;
mem1[2108] = 8'b10010011;
mem1[2109] = 8'b10010011;
mem1[2110] = 8'b10010011;
mem1[2111] = 8'b10010011;
mem1[2112] = 8'b10010100;
mem1[2113] = 8'b10010100;
mem1[2114] = 8'b10010100;
mem1[2115] = 8'b10010100;
mem1[2116] = 8'b10010100;
mem1[2117] = 8'b10010100;
mem1[2118] = 8'b10010100;
mem1[2119] = 8'b10010100;
mem1[2120] = 8'b10010100;
mem1[2121] = 8'b10010101;
mem1[2122] = 8'b10010101;
mem1[2123] = 8'b10010101;
mem1[2124] = 8'b10010101;
mem1[2125] = 8'b10010101;
mem1[2126] = 8'b10010101;
mem1[2127] = 8'b10010101;
mem1[2128] = 8'b10010101;
mem1[2129] = 8'b10010101;
mem1[2130] = 8'b10010101;
mem1[2131] = 8'b10010110;
mem1[2132] = 8'b10010110;
mem1[2133] = 8'b10010110;
mem1[2134] = 8'b10010110;
mem1[2135] = 8'b10010110;
mem1[2136] = 8'b10010110;
mem1[2137] = 8'b10010110;
mem1[2138] = 8'b10010110;
mem1[2139] = 8'b10010110;
mem1[2140] = 8'b10010110;
mem1[2141] = 8'b10010111;
mem1[2142] = 8'b10010111;
mem1[2143] = 8'b10010111;
mem1[2144] = 8'b10010111;
mem1[2145] = 8'b10010111;
mem1[2146] = 8'b10010111;
mem1[2147] = 8'b10010111;
mem1[2148] = 8'b10010111;
mem1[2149] = 8'b10010111;
mem1[2150] = 8'b10010111;
mem1[2151] = 8'b10011000;
mem1[2152] = 8'b10011000;
mem1[2153] = 8'b10011000;
mem1[2154] = 8'b10011000;
mem1[2155] = 8'b10011000;
mem1[2156] = 8'b10011000;
mem1[2157] = 8'b10011000;
mem1[2158] = 8'b10011000;
mem1[2159] = 8'b10011000;
mem1[2160] = 8'b10011001;
mem1[2161] = 8'b10011001;
mem1[2162] = 8'b10011001;
mem1[2163] = 8'b10011001;
mem1[2164] = 8'b10011001;
mem1[2165] = 8'b10011001;
mem1[2166] = 8'b10011001;
mem1[2167] = 8'b10011001;
mem1[2168] = 8'b10011001;
mem1[2169] = 8'b10011001;
mem1[2170] = 8'b10011010;
mem1[2171] = 8'b10011010;
mem1[2172] = 8'b10011010;
mem1[2173] = 8'b10011010;
mem1[2174] = 8'b10011010;
mem1[2175] = 8'b10011010;
mem1[2176] = 8'b10011010;
mem1[2177] = 8'b10011010;
mem1[2178] = 8'b10011010;
mem1[2179] = 8'b10011010;
mem1[2180] = 8'b10011011;
mem1[2181] = 8'b10011011;
mem1[2182] = 8'b10011011;
mem1[2183] = 8'b10011011;
mem1[2184] = 8'b10011011;
mem1[2185] = 8'b10011011;
mem1[2186] = 8'b10011011;
mem1[2187] = 8'b10011011;
mem1[2188] = 8'b10011011;
mem1[2189] = 8'b10011011;
mem1[2190] = 8'b10011100;
mem1[2191] = 8'b10011100;
mem1[2192] = 8'b10011100;
mem1[2193] = 8'b10011100;
mem1[2194] = 8'b10011100;
mem1[2195] = 8'b10011100;
mem1[2196] = 8'b10011100;
mem1[2197] = 8'b10011100;
mem1[2198] = 8'b10011100;
mem1[2199] = 8'b10011101;
mem1[2200] = 8'b10011101;
mem1[2201] = 8'b10011101;
mem1[2202] = 8'b10011101;
mem1[2203] = 8'b10011101;
mem1[2204] = 8'b10011101;
mem1[2205] = 8'b10011101;
mem1[2206] = 8'b10011101;
mem1[2207] = 8'b10011101;
mem1[2208] = 8'b10011101;
mem1[2209] = 8'b10011110;
mem1[2210] = 8'b10011110;
mem1[2211] = 8'b10011110;
mem1[2212] = 8'b10011110;
mem1[2213] = 8'b10011110;
mem1[2214] = 8'b10011110;
mem1[2215] = 8'b10011110;
mem1[2216] = 8'b10011110;
mem1[2217] = 8'b10011110;
mem1[2218] = 8'b10011110;
mem1[2219] = 8'b10011111;
mem1[2220] = 8'b10011111;
mem1[2221] = 8'b10011111;
mem1[2222] = 8'b10011111;
mem1[2223] = 8'b10011111;
mem1[2224] = 8'b10011111;
mem1[2225] = 8'b10011111;
mem1[2226] = 8'b10011111;
mem1[2227] = 8'b10011111;
mem1[2228] = 8'b10011111;
mem1[2229] = 8'b10100000;
mem1[2230] = 8'b10100000;
mem1[2231] = 8'b10100000;
mem1[2232] = 8'b10100000;
mem1[2233] = 8'b10100000;
mem1[2234] = 8'b10100000;
mem1[2235] = 8'b10100000;
mem1[2236] = 8'b10100000;
mem1[2237] = 8'b10100000;
mem1[2238] = 8'b10100000;
mem1[2239] = 8'b10100001;
mem1[2240] = 8'b10100001;
mem1[2241] = 8'b10100001;
mem1[2242] = 8'b10100001;
mem1[2243] = 8'b10100001;
mem1[2244] = 8'b10100001;
mem1[2245] = 8'b10100001;
mem1[2246] = 8'b10100001;
mem1[2247] = 8'b10100001;
mem1[2248] = 8'b10100001;
mem1[2249] = 8'b10100010;
mem1[2250] = 8'b10100010;
mem1[2251] = 8'b10100010;
mem1[2252] = 8'b10100010;
mem1[2253] = 8'b10100010;
mem1[2254] = 8'b10100010;
mem1[2255] = 8'b10100010;
mem1[2256] = 8'b10100010;
mem1[2257] = 8'b10100010;
mem1[2258] = 8'b10100011;
mem1[2259] = 8'b10100011;
mem1[2260] = 8'b10100011;
mem1[2261] = 8'b10100011;
mem1[2262] = 8'b10100011;
mem1[2263] = 8'b10100011;
mem1[2264] = 8'b10100011;
mem1[2265] = 8'b10100011;
mem1[2266] = 8'b10100011;
mem1[2267] = 8'b10100011;
mem1[2268] = 8'b10100100;
mem1[2269] = 8'b10100100;
mem1[2270] = 8'b10100100;
mem1[2271] = 8'b10100100;
mem1[2272] = 8'b10100100;
mem1[2273] = 8'b10100100;
mem1[2274] = 8'b10100100;
mem1[2275] = 8'b10100100;
mem1[2276] = 8'b10100100;
mem1[2277] = 8'b10100100;
mem1[2278] = 8'b10100101;
mem1[2279] = 8'b10100101;
mem1[2280] = 8'b10100101;
mem1[2281] = 8'b10100101;
mem1[2282] = 8'b10100101;
mem1[2283] = 8'b10100101;
mem1[2284] = 8'b10100101;
mem1[2285] = 8'b10100101;
mem1[2286] = 8'b10100101;
mem1[2287] = 8'b10100101;
mem1[2288] = 8'b10100110;
mem1[2289] = 8'b10100110;
mem1[2290] = 8'b10100110;
mem1[2291] = 8'b10100110;
mem1[2292] = 8'b10100110;
mem1[2293] = 8'b10100110;
mem1[2294] = 8'b10100110;
mem1[2295] = 8'b10100110;
mem1[2296] = 8'b10100110;
mem1[2297] = 8'b10100110;
mem1[2298] = 8'b10100111;
mem1[2299] = 8'b10100111;
mem1[2300] = 8'b10100111;
mem1[2301] = 8'b10100111;
mem1[2302] = 8'b10100111;
mem1[2303] = 8'b10100111;
mem1[2304] = 8'b10100111;
mem1[2305] = 8'b10100111;
mem1[2306] = 8'b10100111;
mem1[2307] = 8'b10100111;
mem1[2308] = 8'b10101000;
mem1[2309] = 8'b10101000;
mem1[2310] = 8'b10101000;
mem1[2311] = 8'b10101000;
mem1[2312] = 8'b10101000;
mem1[2313] = 8'b10101000;
mem1[2314] = 8'b10101000;
mem1[2315] = 8'b10101000;
mem1[2316] = 8'b10101000;
mem1[2317] = 8'b10101000;
mem1[2318] = 8'b10101001;
mem1[2319] = 8'b10101001;
mem1[2320] = 8'b10101001;
mem1[2321] = 8'b10101001;
mem1[2322] = 8'b10101001;
mem1[2323] = 8'b10101001;
mem1[2324] = 8'b10101001;
mem1[2325] = 8'b10101001;
mem1[2326] = 8'b10101001;
mem1[2327] = 8'b10101001;
mem1[2328] = 8'b10101001;
mem1[2329] = 8'b10101010;
mem1[2330] = 8'b10101010;
mem1[2331] = 8'b10101010;
mem1[2332] = 8'b10101010;
mem1[2333] = 8'b10101010;
mem1[2334] = 8'b10101010;
mem1[2335] = 8'b10101010;
mem1[2336] = 8'b10101010;
mem1[2337] = 8'b10101010;
mem1[2338] = 8'b10101010;
mem1[2339] = 8'b10101011;
mem1[2340] = 8'b10101011;
mem1[2341] = 8'b10101011;
mem1[2342] = 8'b10101011;
mem1[2343] = 8'b10101011;
mem1[2344] = 8'b10101011;
mem1[2345] = 8'b10101011;
mem1[2346] = 8'b10101011;
mem1[2347] = 8'b10101011;
mem1[2348] = 8'b10101011;
mem1[2349] = 8'b10101100;
mem1[2350] = 8'b10101100;
mem1[2351] = 8'b10101100;
mem1[2352] = 8'b10101100;
mem1[2353] = 8'b10101100;
mem1[2354] = 8'b10101100;
mem1[2355] = 8'b10101100;
mem1[2356] = 8'b10101100;
mem1[2357] = 8'b10101100;
mem1[2358] = 8'b10101100;
mem1[2359] = 8'b10101101;
mem1[2360] = 8'b10101101;
mem1[2361] = 8'b10101101;
mem1[2362] = 8'b10101101;
mem1[2363] = 8'b10101101;
mem1[2364] = 8'b10101101;
mem1[2365] = 8'b10101101;
mem1[2366] = 8'b10101101;
mem1[2367] = 8'b10101101;
mem1[2368] = 8'b10101101;
mem1[2369] = 8'b10101110;
mem1[2370] = 8'b10101110;
mem1[2371] = 8'b10101110;
mem1[2372] = 8'b10101110;
mem1[2373] = 8'b10101110;
mem1[2374] = 8'b10101110;
mem1[2375] = 8'b10101110;
mem1[2376] = 8'b10101110;
mem1[2377] = 8'b10101110;
mem1[2378] = 8'b10101110;
mem1[2379] = 8'b10101110;
mem1[2380] = 8'b10101111;
mem1[2381] = 8'b10101111;
mem1[2382] = 8'b10101111;
mem1[2383] = 8'b10101111;
mem1[2384] = 8'b10101111;
mem1[2385] = 8'b10101111;
mem1[2386] = 8'b10101111;
mem1[2387] = 8'b10101111;
mem1[2388] = 8'b10101111;
mem1[2389] = 8'b10101111;
mem1[2390] = 8'b10110000;
mem1[2391] = 8'b10110000;
mem1[2392] = 8'b10110000;
mem1[2393] = 8'b10110000;
mem1[2394] = 8'b10110000;
mem1[2395] = 8'b10110000;
mem1[2396] = 8'b10110000;
mem1[2397] = 8'b10110000;
mem1[2398] = 8'b10110000;
mem1[2399] = 8'b10110000;
mem1[2400] = 8'b10110001;
mem1[2401] = 8'b10110001;
mem1[2402] = 8'b10110001;
mem1[2403] = 8'b10110001;
mem1[2404] = 8'b10110001;
mem1[2405] = 8'b10110001;
mem1[2406] = 8'b10110001;
mem1[2407] = 8'b10110001;
mem1[2408] = 8'b10110001;
mem1[2409] = 8'b10110001;
mem1[2410] = 8'b10110010;
mem1[2411] = 8'b10110010;
mem1[2412] = 8'b10110010;
mem1[2413] = 8'b10110010;
mem1[2414] = 8'b10110010;
mem1[2415] = 8'b10110010;
mem1[2416] = 8'b10110010;
mem1[2417] = 8'b10110010;
mem1[2418] = 8'b10110010;
mem1[2419] = 8'b10110010;
mem1[2420] = 8'b10110010;
mem1[2421] = 8'b10110011;
mem1[2422] = 8'b10110011;
mem1[2423] = 8'b10110011;
mem1[2424] = 8'b10110011;
mem1[2425] = 8'b10110011;
mem1[2426] = 8'b10110011;
mem1[2427] = 8'b10110011;
mem1[2428] = 8'b10110011;
mem1[2429] = 8'b10110011;
mem1[2430] = 8'b10110011;
mem1[2431] = 8'b10110100;
mem1[2432] = 8'b10110100;
mem1[2433] = 8'b10110100;
mem1[2434] = 8'b10110100;
mem1[2435] = 8'b10110100;
mem1[2436] = 8'b10110100;
mem1[2437] = 8'b10110100;
mem1[2438] = 8'b10110100;
mem1[2439] = 8'b10110100;
mem1[2440] = 8'b10110100;
mem1[2441] = 8'b10110100;
mem1[2442] = 8'b10110101;
mem1[2443] = 8'b10110101;
mem1[2444] = 8'b10110101;
mem1[2445] = 8'b10110101;
mem1[2446] = 8'b10110101;
mem1[2447] = 8'b10110101;
mem1[2448] = 8'b10110101;
mem1[2449] = 8'b10110101;
mem1[2450] = 8'b10110101;
mem1[2451] = 8'b10110101;
mem1[2452] = 8'b10110110;
mem1[2453] = 8'b10110110;
mem1[2454] = 8'b10110110;
mem1[2455] = 8'b10110110;
mem1[2456] = 8'b10110110;
mem1[2457] = 8'b10110110;
mem1[2458] = 8'b10110110;
mem1[2459] = 8'b10110110;
mem1[2460] = 8'b10110110;
mem1[2461] = 8'b10110110;
mem1[2462] = 8'b10110110;
mem1[2463] = 8'b10110111;
mem1[2464] = 8'b10110111;
mem1[2465] = 8'b10110111;
mem1[2466] = 8'b10110111;
mem1[2467] = 8'b10110111;
mem1[2468] = 8'b10110111;
mem1[2469] = 8'b10110111;
mem1[2470] = 8'b10110111;
mem1[2471] = 8'b10110111;
mem1[2472] = 8'b10110111;
mem1[2473] = 8'b10111000;
mem1[2474] = 8'b10111000;
mem1[2475] = 8'b10111000;
mem1[2476] = 8'b10111000;
mem1[2477] = 8'b10111000;
mem1[2478] = 8'b10111000;
mem1[2479] = 8'b10111000;
mem1[2480] = 8'b10111000;
mem1[2481] = 8'b10111000;
mem1[2482] = 8'b10111000;
mem1[2483] = 8'b10111000;
mem1[2484] = 8'b10111001;
mem1[2485] = 8'b10111001;
mem1[2486] = 8'b10111001;
mem1[2487] = 8'b10111001;
mem1[2488] = 8'b10111001;
mem1[2489] = 8'b10111001;
mem1[2490] = 8'b10111001;
mem1[2491] = 8'b10111001;
mem1[2492] = 8'b10111001;
mem1[2493] = 8'b10111001;
mem1[2494] = 8'b10111001;
mem1[2495] = 8'b10111010;
mem1[2496] = 8'b10111010;
mem1[2497] = 8'b10111010;
mem1[2498] = 8'b10111010;
mem1[2499] = 8'b10111010;
mem1[2500] = 8'b10111010;
mem1[2501] = 8'b10111010;
mem1[2502] = 8'b10111010;
mem1[2503] = 8'b10111010;
mem1[2504] = 8'b10111010;
mem1[2505] = 8'b10111011;
mem1[2506] = 8'b10111011;
mem1[2507] = 8'b10111011;
mem1[2508] = 8'b10111011;
mem1[2509] = 8'b10111011;
mem1[2510] = 8'b10111011;
mem1[2511] = 8'b10111011;
mem1[2512] = 8'b10111011;
mem1[2513] = 8'b10111011;
mem1[2514] = 8'b10111011;
mem1[2515] = 8'b10111011;
mem1[2516] = 8'b10111100;
mem1[2517] = 8'b10111100;
mem1[2518] = 8'b10111100;
mem1[2519] = 8'b10111100;
mem1[2520] = 8'b10111100;
mem1[2521] = 8'b10111100;
mem1[2522] = 8'b10111100;
mem1[2523] = 8'b10111100;
mem1[2524] = 8'b10111100;
mem1[2525] = 8'b10111100;
mem1[2526] = 8'b10111100;
mem1[2527] = 8'b10111101;
mem1[2528] = 8'b10111101;
mem1[2529] = 8'b10111101;
mem1[2530] = 8'b10111101;
mem1[2531] = 8'b10111101;
mem1[2532] = 8'b10111101;
mem1[2533] = 8'b10111101;
mem1[2534] = 8'b10111101;
mem1[2535] = 8'b10111101;
mem1[2536] = 8'b10111101;
mem1[2537] = 8'b10111101;
mem1[2538] = 8'b10111110;
mem1[2539] = 8'b10111110;
mem1[2540] = 8'b10111110;
mem1[2541] = 8'b10111110;
mem1[2542] = 8'b10111110;
mem1[2543] = 8'b10111110;
mem1[2544] = 8'b10111110;
mem1[2545] = 8'b10111110;
mem1[2546] = 8'b10111110;
mem1[2547] = 8'b10111110;
mem1[2548] = 8'b10111110;
mem1[2549] = 8'b10111111;
mem1[2550] = 8'b10111111;
mem1[2551] = 8'b10111111;
mem1[2552] = 8'b10111111;
mem1[2553] = 8'b10111111;
mem1[2554] = 8'b10111111;
mem1[2555] = 8'b10111111;
mem1[2556] = 8'b10111111;
mem1[2557] = 8'b10111111;
mem1[2558] = 8'b10111111;
mem1[2559] = 8'b10111111;
mem1[2560] = 8'b11000000;
mem1[2561] = 8'b11000000;
mem1[2562] = 8'b11000000;
mem1[2563] = 8'b11000000;
mem1[2564] = 8'b11000000;
mem1[2565] = 8'b11000000;
mem1[2566] = 8'b11000000;
mem1[2567] = 8'b11000000;
mem1[2568] = 8'b11000000;
mem1[2569] = 8'b11000000;
mem1[2570] = 8'b11000000;
mem1[2571] = 8'b11000001;
mem1[2572] = 8'b11000001;
mem1[2573] = 8'b11000001;
mem1[2574] = 8'b11000001;
mem1[2575] = 8'b11000001;
mem1[2576] = 8'b11000001;
mem1[2577] = 8'b11000001;
mem1[2578] = 8'b11000001;
mem1[2579] = 8'b11000001;
mem1[2580] = 8'b11000001;
mem1[2581] = 8'b11000001;
mem1[2582] = 8'b11000010;
mem1[2583] = 8'b11000010;
mem1[2584] = 8'b11000010;
mem1[2585] = 8'b11000010;
mem1[2586] = 8'b11000010;
mem1[2587] = 8'b11000010;
mem1[2588] = 8'b11000010;
mem1[2589] = 8'b11000010;
mem1[2590] = 8'b11000010;
mem1[2591] = 8'b11000010;
mem1[2592] = 8'b11000010;
mem1[2593] = 8'b11000011;
mem1[2594] = 8'b11000011;
mem1[2595] = 8'b11000011;
mem1[2596] = 8'b11000011;
mem1[2597] = 8'b11000011;
mem1[2598] = 8'b11000011;
mem1[2599] = 8'b11000011;
mem1[2600] = 8'b11000011;
mem1[2601] = 8'b11000011;
mem1[2602] = 8'b11000011;
mem1[2603] = 8'b11000011;
mem1[2604] = 8'b11000100;
mem1[2605] = 8'b11000100;
mem1[2606] = 8'b11000100;
mem1[2607] = 8'b11000100;
mem1[2608] = 8'b11000100;
mem1[2609] = 8'b11000100;
mem1[2610] = 8'b11000100;
mem1[2611] = 8'b11000100;
mem1[2612] = 8'b11000100;
mem1[2613] = 8'b11000100;
mem1[2614] = 8'b11000100;
mem1[2615] = 8'b11000100;
mem1[2616] = 8'b11000101;
mem1[2617] = 8'b11000101;
mem1[2618] = 8'b11000101;
mem1[2619] = 8'b11000101;
mem1[2620] = 8'b11000101;
mem1[2621] = 8'b11000101;
mem1[2622] = 8'b11000101;
mem1[2623] = 8'b11000101;
mem1[2624] = 8'b11000101;
mem1[2625] = 8'b11000101;
mem1[2626] = 8'b11000101;
mem1[2627] = 8'b11000110;
mem1[2628] = 8'b11000110;
mem1[2629] = 8'b11000110;
mem1[2630] = 8'b11000110;
mem1[2631] = 8'b11000110;
mem1[2632] = 8'b11000110;
mem1[2633] = 8'b11000110;
mem1[2634] = 8'b11000110;
mem1[2635] = 8'b11000110;
mem1[2636] = 8'b11000110;
mem1[2637] = 8'b11000110;
mem1[2638] = 8'b11000110;
mem1[2639] = 8'b11000111;
mem1[2640] = 8'b11000111;
mem1[2641] = 8'b11000111;
mem1[2642] = 8'b11000111;
mem1[2643] = 8'b11000111;
mem1[2644] = 8'b11000111;
mem1[2645] = 8'b11000111;
mem1[2646] = 8'b11000111;
mem1[2647] = 8'b11000111;
mem1[2648] = 8'b11000111;
mem1[2649] = 8'b11000111;
mem1[2650] = 8'b11001000;
mem1[2651] = 8'b11001000;
mem1[2652] = 8'b11001000;
mem1[2653] = 8'b11001000;
mem1[2654] = 8'b11001000;
mem1[2655] = 8'b11001000;
mem1[2656] = 8'b11001000;
mem1[2657] = 8'b11001000;
mem1[2658] = 8'b11001000;
mem1[2659] = 8'b11001000;
mem1[2660] = 8'b11001000;
mem1[2661] = 8'b11001000;
mem1[2662] = 8'b11001001;
mem1[2663] = 8'b11001001;
mem1[2664] = 8'b11001001;
mem1[2665] = 8'b11001001;
mem1[2666] = 8'b11001001;
mem1[2667] = 8'b11001001;
mem1[2668] = 8'b11001001;
mem1[2669] = 8'b11001001;
mem1[2670] = 8'b11001001;
mem1[2671] = 8'b11001001;
mem1[2672] = 8'b11001001;
mem1[2673] = 8'b11001010;
mem1[2674] = 8'b11001010;
mem1[2675] = 8'b11001010;
mem1[2676] = 8'b11001010;
mem1[2677] = 8'b11001010;
mem1[2678] = 8'b11001010;
mem1[2679] = 8'b11001010;
mem1[2680] = 8'b11001010;
mem1[2681] = 8'b11001010;
mem1[2682] = 8'b11001010;
mem1[2683] = 8'b11001010;
mem1[2684] = 8'b11001010;
mem1[2685] = 8'b11001011;
mem1[2686] = 8'b11001011;
mem1[2687] = 8'b11001011;
mem1[2688] = 8'b11001011;
mem1[2689] = 8'b11001011;
mem1[2690] = 8'b11001011;
mem1[2691] = 8'b11001011;
mem1[2692] = 8'b11001011;
mem1[2693] = 8'b11001011;
mem1[2694] = 8'b11001011;
mem1[2695] = 8'b11001011;
mem1[2696] = 8'b11001011;
mem1[2697] = 8'b11001100;
mem1[2698] = 8'b11001100;
mem1[2699] = 8'b11001100;
mem1[2700] = 8'b11001100;
mem1[2701] = 8'b11001100;
mem1[2702] = 8'b11001100;
mem1[2703] = 8'b11001100;
mem1[2704] = 8'b11001100;
mem1[2705] = 8'b11001100;
mem1[2706] = 8'b11001100;
mem1[2707] = 8'b11001100;
mem1[2708] = 8'b11001100;
mem1[2709] = 8'b11001101;
mem1[2710] = 8'b11001101;
mem1[2711] = 8'b11001101;
mem1[2712] = 8'b11001101;
mem1[2713] = 8'b11001101;
mem1[2714] = 8'b11001101;
mem1[2715] = 8'b11001101;
mem1[2716] = 8'b11001101;
mem1[2717] = 8'b11001101;
mem1[2718] = 8'b11001101;
mem1[2719] = 8'b11001101;
mem1[2720] = 8'b11001101;
mem1[2721] = 8'b11001110;
mem1[2722] = 8'b11001110;
mem1[2723] = 8'b11001110;
mem1[2724] = 8'b11001110;
mem1[2725] = 8'b11001110;
mem1[2726] = 8'b11001110;
mem1[2727] = 8'b11001110;
mem1[2728] = 8'b11001110;
mem1[2729] = 8'b11001110;
mem1[2730] = 8'b11001110;
mem1[2731] = 8'b11001110;
mem1[2732] = 8'b11001110;
mem1[2733] = 8'b11001111;
mem1[2734] = 8'b11001111;
mem1[2735] = 8'b11001111;
mem1[2736] = 8'b11001111;
mem1[2737] = 8'b11001111;
mem1[2738] = 8'b11001111;
mem1[2739] = 8'b11001111;
mem1[2740] = 8'b11001111;
mem1[2741] = 8'b11001111;
mem1[2742] = 8'b11001111;
mem1[2743] = 8'b11001111;
mem1[2744] = 8'b11001111;
mem1[2745] = 8'b11010000;
mem1[2746] = 8'b11010000;
mem1[2747] = 8'b11010000;
mem1[2748] = 8'b11010000;
mem1[2749] = 8'b11010000;
mem1[2750] = 8'b11010000;
mem1[2751] = 8'b11010000;
mem1[2752] = 8'b11010000;
mem1[2753] = 8'b11010000;
mem1[2754] = 8'b11010000;
mem1[2755] = 8'b11010000;
mem1[2756] = 8'b11010000;
mem1[2757] = 8'b11010001;
mem1[2758] = 8'b11010001;
mem1[2759] = 8'b11010001;
mem1[2760] = 8'b11010001;
mem1[2761] = 8'b11010001;
mem1[2762] = 8'b11010001;
mem1[2763] = 8'b11010001;
mem1[2764] = 8'b11010001;
mem1[2765] = 8'b11010001;
mem1[2766] = 8'b11010001;
mem1[2767] = 8'b11010001;
mem1[2768] = 8'b11010001;
mem1[2769] = 8'b11010001;
mem1[2770] = 8'b11010010;
mem1[2771] = 8'b11010010;
mem1[2772] = 8'b11010010;
mem1[2773] = 8'b11010010;
mem1[2774] = 8'b11010010;
mem1[2775] = 8'b11010010;
mem1[2776] = 8'b11010010;
mem1[2777] = 8'b11010010;
mem1[2778] = 8'b11010010;
mem1[2779] = 8'b11010010;
mem1[2780] = 8'b11010010;
mem1[2781] = 8'b11010010;
mem1[2782] = 8'b11010011;
mem1[2783] = 8'b11010011;
mem1[2784] = 8'b11010011;
mem1[2785] = 8'b11010011;
mem1[2786] = 8'b11010011;
mem1[2787] = 8'b11010011;
mem1[2788] = 8'b11010011;
mem1[2789] = 8'b11010011;
mem1[2790] = 8'b11010011;
mem1[2791] = 8'b11010011;
mem1[2792] = 8'b11010011;
mem1[2793] = 8'b11010011;
mem1[2794] = 8'b11010011;
mem1[2795] = 8'b11010100;
mem1[2796] = 8'b11010100;
mem1[2797] = 8'b11010100;
mem1[2798] = 8'b11010100;
mem1[2799] = 8'b11010100;
mem1[2800] = 8'b11010100;
mem1[2801] = 8'b11010100;
mem1[2802] = 8'b11010100;
mem1[2803] = 8'b11010100;
mem1[2804] = 8'b11010100;
mem1[2805] = 8'b11010100;
mem1[2806] = 8'b11010100;
mem1[2807] = 8'b11010100;
mem1[2808] = 8'b11010101;
mem1[2809] = 8'b11010101;
mem1[2810] = 8'b11010101;
mem1[2811] = 8'b11010101;
mem1[2812] = 8'b11010101;
mem1[2813] = 8'b11010101;
mem1[2814] = 8'b11010101;
mem1[2815] = 8'b11010101;
mem1[2816] = 8'b11010101;
mem1[2817] = 8'b11010101;
mem1[2818] = 8'b11010101;
mem1[2819] = 8'b11010101;
mem1[2820] = 8'b11010110;
mem1[2821] = 8'b11010110;
mem1[2822] = 8'b11010110;
mem1[2823] = 8'b11010110;
mem1[2824] = 8'b11010110;
mem1[2825] = 8'b11010110;
mem1[2826] = 8'b11010110;
mem1[2827] = 8'b11010110;
mem1[2828] = 8'b11010110;
mem1[2829] = 8'b11010110;
mem1[2830] = 8'b11010110;
mem1[2831] = 8'b11010110;
mem1[2832] = 8'b11010110;
mem1[2833] = 8'b11010111;
mem1[2834] = 8'b11010111;
mem1[2835] = 8'b11010111;
mem1[2836] = 8'b11010111;
mem1[2837] = 8'b11010111;
mem1[2838] = 8'b11010111;
mem1[2839] = 8'b11010111;
mem1[2840] = 8'b11010111;
mem1[2841] = 8'b11010111;
mem1[2842] = 8'b11010111;
mem1[2843] = 8'b11010111;
mem1[2844] = 8'b11010111;
mem1[2845] = 8'b11010111;
mem1[2846] = 8'b11011000;
mem1[2847] = 8'b11011000;
mem1[2848] = 8'b11011000;
mem1[2849] = 8'b11011000;
mem1[2850] = 8'b11011000;
mem1[2851] = 8'b11011000;
mem1[2852] = 8'b11011000;
mem1[2853] = 8'b11011000;
mem1[2854] = 8'b11011000;
mem1[2855] = 8'b11011000;
mem1[2856] = 8'b11011000;
mem1[2857] = 8'b11011000;
mem1[2858] = 8'b11011000;
mem1[2859] = 8'b11011000;
mem1[2860] = 8'b11011001;
mem1[2861] = 8'b11011001;
mem1[2862] = 8'b11011001;
mem1[2863] = 8'b11011001;
mem1[2864] = 8'b11011001;
mem1[2865] = 8'b11011001;
mem1[2866] = 8'b11011001;
mem1[2867] = 8'b11011001;
mem1[2868] = 8'b11011001;
mem1[2869] = 8'b11011001;
mem1[2870] = 8'b11011001;
mem1[2871] = 8'b11011001;
mem1[2872] = 8'b11011001;
mem1[2873] = 8'b11011010;
mem1[2874] = 8'b11011010;
mem1[2875] = 8'b11011010;
mem1[2876] = 8'b11011010;
mem1[2877] = 8'b11011010;
mem1[2878] = 8'b11011010;
mem1[2879] = 8'b11011010;
mem1[2880] = 8'b11011010;
mem1[2881] = 8'b11011010;
mem1[2882] = 8'b11011010;
mem1[2883] = 8'b11011010;
mem1[2884] = 8'b11011010;
mem1[2885] = 8'b11011010;
mem1[2886] = 8'b11011010;
mem1[2887] = 8'b11011011;
mem1[2888] = 8'b11011011;
mem1[2889] = 8'b11011011;
mem1[2890] = 8'b11011011;
mem1[2891] = 8'b11011011;
mem1[2892] = 8'b11011011;
mem1[2893] = 8'b11011011;
mem1[2894] = 8'b11011011;
mem1[2895] = 8'b11011011;
mem1[2896] = 8'b11011011;
mem1[2897] = 8'b11011011;
mem1[2898] = 8'b11011011;
mem1[2899] = 8'b11011011;
mem1[2900] = 8'b11011100;
mem1[2901] = 8'b11011100;
mem1[2902] = 8'b11011100;
mem1[2903] = 8'b11011100;
mem1[2904] = 8'b11011100;
mem1[2905] = 8'b11011100;
mem1[2906] = 8'b11011100;
mem1[2907] = 8'b11011100;
mem1[2908] = 8'b11011100;
mem1[2909] = 8'b11011100;
mem1[2910] = 8'b11011100;
mem1[2911] = 8'b11011100;
mem1[2912] = 8'b11011100;
mem1[2913] = 8'b11011100;
mem1[2914] = 8'b11011101;
mem1[2915] = 8'b11011101;
mem1[2916] = 8'b11011101;
mem1[2917] = 8'b11011101;
mem1[2918] = 8'b11011101;
mem1[2919] = 8'b11011101;
mem1[2920] = 8'b11011101;
mem1[2921] = 8'b11011101;
mem1[2922] = 8'b11011101;
mem1[2923] = 8'b11011101;
mem1[2924] = 8'b11011101;
mem1[2925] = 8'b11011101;
mem1[2926] = 8'b11011101;
mem1[2927] = 8'b11011101;
mem1[2928] = 8'b11011110;
mem1[2929] = 8'b11011110;
mem1[2930] = 8'b11011110;
mem1[2931] = 8'b11011110;
mem1[2932] = 8'b11011110;
mem1[2933] = 8'b11011110;
mem1[2934] = 8'b11011110;
mem1[2935] = 8'b11011110;
mem1[2936] = 8'b11011110;
mem1[2937] = 8'b11011110;
mem1[2938] = 8'b11011110;
mem1[2939] = 8'b11011110;
mem1[2940] = 8'b11011110;
mem1[2941] = 8'b11011110;
mem1[2942] = 8'b11011111;
mem1[2943] = 8'b11011111;
mem1[2944] = 8'b11011111;
mem1[2945] = 8'b11011111;
mem1[2946] = 8'b11011111;
mem1[2947] = 8'b11011111;
mem1[2948] = 8'b11011111;
mem1[2949] = 8'b11011111;
mem1[2950] = 8'b11011111;
mem1[2951] = 8'b11011111;
mem1[2952] = 8'b11011111;
mem1[2953] = 8'b11011111;
mem1[2954] = 8'b11011111;
mem1[2955] = 8'b11011111;
mem1[2956] = 8'b11100000;
mem1[2957] = 8'b11100000;
mem1[2958] = 8'b11100000;
mem1[2959] = 8'b11100000;
mem1[2960] = 8'b11100000;
mem1[2961] = 8'b11100000;
mem1[2962] = 8'b11100000;
mem1[2963] = 8'b11100000;
mem1[2964] = 8'b11100000;
mem1[2965] = 8'b11100000;
mem1[2966] = 8'b11100000;
mem1[2967] = 8'b11100000;
mem1[2968] = 8'b11100000;
mem1[2969] = 8'b11100000;
mem1[2970] = 8'b11100000;
mem1[2971] = 8'b11100001;
mem1[2972] = 8'b11100001;
mem1[2973] = 8'b11100001;
mem1[2974] = 8'b11100001;
mem1[2975] = 8'b11100001;
mem1[2976] = 8'b11100001;
mem1[2977] = 8'b11100001;
mem1[2978] = 8'b11100001;
mem1[2979] = 8'b11100001;
mem1[2980] = 8'b11100001;
mem1[2981] = 8'b11100001;
mem1[2982] = 8'b11100001;
mem1[2983] = 8'b11100001;
mem1[2984] = 8'b11100001;
mem1[2985] = 8'b11100001;
mem1[2986] = 8'b11100010;
mem1[2987] = 8'b11100010;
mem1[2988] = 8'b11100010;
mem1[2989] = 8'b11100010;
mem1[2990] = 8'b11100010;
mem1[2991] = 8'b11100010;
mem1[2992] = 8'b11100010;
mem1[2993] = 8'b11100010;
mem1[2994] = 8'b11100010;
mem1[2995] = 8'b11100010;
mem1[2996] = 8'b11100010;
mem1[2997] = 8'b11100010;
mem1[2998] = 8'b11100010;
mem1[2999] = 8'b11100010;
mem1[3000] = 8'b11100010;
mem1[3001] = 8'b11100011;
mem1[3002] = 8'b11100011;
mem1[3003] = 8'b11100011;
mem1[3004] = 8'b11100011;
mem1[3005] = 8'b11100011;
mem1[3006] = 8'b11100011;
mem1[3007] = 8'b11100011;
mem1[3008] = 8'b11100011;
mem1[3009] = 8'b11100011;
mem1[3010] = 8'b11100011;
mem1[3011] = 8'b11100011;
mem1[3012] = 8'b11100011;
mem1[3013] = 8'b11100011;
mem1[3014] = 8'b11100011;
mem1[3015] = 8'b11100011;
mem1[3016] = 8'b11100100;
mem1[3017] = 8'b11100100;
mem1[3018] = 8'b11100100;
mem1[3019] = 8'b11100100;
mem1[3020] = 8'b11100100;
mem1[3021] = 8'b11100100;
mem1[3022] = 8'b11100100;
mem1[3023] = 8'b11100100;
mem1[3024] = 8'b11100100;
mem1[3025] = 8'b11100100;
mem1[3026] = 8'b11100100;
mem1[3027] = 8'b11100100;
mem1[3028] = 8'b11100100;
mem1[3029] = 8'b11100100;
mem1[3030] = 8'b11100100;
mem1[3031] = 8'b11100101;
mem1[3032] = 8'b11100101;
mem1[3033] = 8'b11100101;
mem1[3034] = 8'b11100101;
mem1[3035] = 8'b11100101;
mem1[3036] = 8'b11100101;
mem1[3037] = 8'b11100101;
mem1[3038] = 8'b11100101;
mem1[3039] = 8'b11100101;
mem1[3040] = 8'b11100101;
mem1[3041] = 8'b11100101;
mem1[3042] = 8'b11100101;
mem1[3043] = 8'b11100101;
mem1[3044] = 8'b11100101;
mem1[3045] = 8'b11100101;
mem1[3046] = 8'b11100101;
mem1[3047] = 8'b11100110;
mem1[3048] = 8'b11100110;
mem1[3049] = 8'b11100110;
mem1[3050] = 8'b11100110;
mem1[3051] = 8'b11100110;
mem1[3052] = 8'b11100110;
mem1[3053] = 8'b11100110;
mem1[3054] = 8'b11100110;
mem1[3055] = 8'b11100110;
mem1[3056] = 8'b11100110;
mem1[3057] = 8'b11100110;
mem1[3058] = 8'b11100110;
mem1[3059] = 8'b11100110;
mem1[3060] = 8'b11100110;
mem1[3061] = 8'b11100110;
mem1[3062] = 8'b11100110;
mem1[3063] = 8'b11100111;
mem1[3064] = 8'b11100111;
mem1[3065] = 8'b11100111;
mem1[3066] = 8'b11100111;
mem1[3067] = 8'b11100111;
mem1[3068] = 8'b11100111;
mem1[3069] = 8'b11100111;
mem1[3070] = 8'b11100111;
mem1[3071] = 8'b11100111;
mem1[3072] = 8'b11100111;
mem1[3073] = 8'b11100111;
mem1[3074] = 8'b11100111;
mem1[3075] = 8'b11100111;
mem1[3076] = 8'b11100111;
mem1[3077] = 8'b11100111;
mem1[3078] = 8'b11100111;
mem1[3079] = 8'b11101000;
mem1[3080] = 8'b11101000;
mem1[3081] = 8'b11101000;
mem1[3082] = 8'b11101000;
mem1[3083] = 8'b11101000;
mem1[3084] = 8'b11101000;
mem1[3085] = 8'b11101000;
mem1[3086] = 8'b11101000;
mem1[3087] = 8'b11101000;
mem1[3088] = 8'b11101000;
mem1[3089] = 8'b11101000;
mem1[3090] = 8'b11101000;
mem1[3091] = 8'b11101000;
mem1[3092] = 8'b11101000;
mem1[3093] = 8'b11101000;
mem1[3094] = 8'b11101000;
mem1[3095] = 8'b11101000;
mem1[3096] = 8'b11101001;
mem1[3097] = 8'b11101001;
mem1[3098] = 8'b11101001;
mem1[3099] = 8'b11101001;
mem1[3100] = 8'b11101001;
mem1[3101] = 8'b11101001;
mem1[3102] = 8'b11101001;
mem1[3103] = 8'b11101001;
mem1[3104] = 8'b11101001;
mem1[3105] = 8'b11101001;
mem1[3106] = 8'b11101001;
mem1[3107] = 8'b11101001;
mem1[3108] = 8'b11101001;
mem1[3109] = 8'b11101001;
mem1[3110] = 8'b11101001;
mem1[3111] = 8'b11101001;
mem1[3112] = 8'b11101001;
mem1[3113] = 8'b11101010;
mem1[3114] = 8'b11101010;
mem1[3115] = 8'b11101010;
mem1[3116] = 8'b11101010;
mem1[3117] = 8'b11101010;
mem1[3118] = 8'b11101010;
mem1[3119] = 8'b11101010;
mem1[3120] = 8'b11101010;
mem1[3121] = 8'b11101010;
mem1[3122] = 8'b11101010;
mem1[3123] = 8'b11101010;
mem1[3124] = 8'b11101010;
mem1[3125] = 8'b11101010;
mem1[3126] = 8'b11101010;
mem1[3127] = 8'b11101010;
mem1[3128] = 8'b11101010;
mem1[3129] = 8'b11101010;
mem1[3130] = 8'b11101011;
mem1[3131] = 8'b11101011;
mem1[3132] = 8'b11101011;
mem1[3133] = 8'b11101011;
mem1[3134] = 8'b11101011;
mem1[3135] = 8'b11101011;
mem1[3136] = 8'b11101011;
mem1[3137] = 8'b11101011;
mem1[3138] = 8'b11101011;
mem1[3139] = 8'b11101011;
mem1[3140] = 8'b11101011;
mem1[3141] = 8'b11101011;
mem1[3142] = 8'b11101011;
mem1[3143] = 8'b11101011;
mem1[3144] = 8'b11101011;
mem1[3145] = 8'b11101011;
mem1[3146] = 8'b11101011;
mem1[3147] = 8'b11101100;
mem1[3148] = 8'b11101100;
mem1[3149] = 8'b11101100;
mem1[3150] = 8'b11101100;
mem1[3151] = 8'b11101100;
mem1[3152] = 8'b11101100;
mem1[3153] = 8'b11101100;
mem1[3154] = 8'b11101100;
mem1[3155] = 8'b11101100;
mem1[3156] = 8'b11101100;
mem1[3157] = 8'b11101100;
mem1[3158] = 8'b11101100;
mem1[3159] = 8'b11101100;
mem1[3160] = 8'b11101100;
mem1[3161] = 8'b11101100;
mem1[3162] = 8'b11101100;
mem1[3163] = 8'b11101100;
mem1[3164] = 8'b11101100;
mem1[3165] = 8'b11101101;
mem1[3166] = 8'b11101101;
mem1[3167] = 8'b11101101;
mem1[3168] = 8'b11101101;
mem1[3169] = 8'b11101101;
mem1[3170] = 8'b11101101;
mem1[3171] = 8'b11101101;
mem1[3172] = 8'b11101101;
mem1[3173] = 8'b11101101;
mem1[3174] = 8'b11101101;
mem1[3175] = 8'b11101101;
mem1[3176] = 8'b11101101;
mem1[3177] = 8'b11101101;
mem1[3178] = 8'b11101101;
mem1[3179] = 8'b11101101;
mem1[3180] = 8'b11101101;
mem1[3181] = 8'b11101101;
mem1[3182] = 8'b11101101;
mem1[3183] = 8'b11101101;
mem1[3184] = 8'b11101110;
mem1[3185] = 8'b11101110;
mem1[3186] = 8'b11101110;
mem1[3187] = 8'b11101110;
mem1[3188] = 8'b11101110;
mem1[3189] = 8'b11101110;
mem1[3190] = 8'b11101110;
mem1[3191] = 8'b11101110;
mem1[3192] = 8'b11101110;
mem1[3193] = 8'b11101110;
mem1[3194] = 8'b11101110;
mem1[3195] = 8'b11101110;
mem1[3196] = 8'b11101110;
mem1[3197] = 8'b11101110;
mem1[3198] = 8'b11101110;
mem1[3199] = 8'b11101110;
mem1[3200] = 8'b11101110;
mem1[3201] = 8'b11101110;
mem1[3202] = 8'b11101110;
mem1[3203] = 8'b11101111;
mem1[3204] = 8'b11101111;
mem1[3205] = 8'b11101111;
mem1[3206] = 8'b11101111;
mem1[3207] = 8'b11101111;
mem1[3208] = 8'b11101111;
mem1[3209] = 8'b11101111;
mem1[3210] = 8'b11101111;
mem1[3211] = 8'b11101111;
mem1[3212] = 8'b11101111;
mem1[3213] = 8'b11101111;
mem1[3214] = 8'b11101111;
mem1[3215] = 8'b11101111;
mem1[3216] = 8'b11101111;
mem1[3217] = 8'b11101111;
mem1[3218] = 8'b11101111;
mem1[3219] = 8'b11101111;
mem1[3220] = 8'b11101111;
mem1[3221] = 8'b11101111;
mem1[3222] = 8'b11110000;
mem1[3223] = 8'b11110000;
mem1[3224] = 8'b11110000;
mem1[3225] = 8'b11110000;
mem1[3226] = 8'b11110000;
mem1[3227] = 8'b11110000;
mem1[3228] = 8'b11110000;
mem1[3229] = 8'b11110000;
mem1[3230] = 8'b11110000;
mem1[3231] = 8'b11110000;
mem1[3232] = 8'b11110000;
mem1[3233] = 8'b11110000;
mem1[3234] = 8'b11110000;
mem1[3235] = 8'b11110000;
mem1[3236] = 8'b11110000;
mem1[3237] = 8'b11110000;
mem1[3238] = 8'b11110000;
mem1[3239] = 8'b11110000;
mem1[3240] = 8'b11110000;
mem1[3241] = 8'b11110000;
mem1[3242] = 8'b11110001;
mem1[3243] = 8'b11110001;
mem1[3244] = 8'b11110001;
mem1[3245] = 8'b11110001;
mem1[3246] = 8'b11110001;
mem1[3247] = 8'b11110001;
mem1[3248] = 8'b11110001;
mem1[3249] = 8'b11110001;
mem1[3250] = 8'b11110001;
mem1[3251] = 8'b11110001;
mem1[3252] = 8'b11110001;
mem1[3253] = 8'b11110001;
mem1[3254] = 8'b11110001;
mem1[3255] = 8'b11110001;
mem1[3256] = 8'b11110001;
mem1[3257] = 8'b11110001;
mem1[3258] = 8'b11110001;
mem1[3259] = 8'b11110001;
mem1[3260] = 8'b11110001;
mem1[3261] = 8'b11110001;
mem1[3262] = 8'b11110001;
mem1[3263] = 8'b11110010;
mem1[3264] = 8'b11110010;
mem1[3265] = 8'b11110010;
mem1[3266] = 8'b11110010;
mem1[3267] = 8'b11110010;
mem1[3268] = 8'b11110010;
mem1[3269] = 8'b11110010;
mem1[3270] = 8'b11110010;
mem1[3271] = 8'b11110010;
mem1[3272] = 8'b11110010;
mem1[3273] = 8'b11110010;
mem1[3274] = 8'b11110010;
mem1[3275] = 8'b11110010;
mem1[3276] = 8'b11110010;
mem1[3277] = 8'b11110010;
mem1[3278] = 8'b11110010;
mem1[3279] = 8'b11110010;
mem1[3280] = 8'b11110010;
mem1[3281] = 8'b11110010;
mem1[3282] = 8'b11110010;
mem1[3283] = 8'b11110010;
mem1[3284] = 8'b11110011;
mem1[3285] = 8'b11110011;
mem1[3286] = 8'b11110011;
mem1[3287] = 8'b11110011;
mem1[3288] = 8'b11110011;
mem1[3289] = 8'b11110011;
mem1[3290] = 8'b11110011;
mem1[3291] = 8'b11110011;
mem1[3292] = 8'b11110011;
mem1[3293] = 8'b11110011;
mem1[3294] = 8'b11110011;
mem1[3295] = 8'b11110011;
mem1[3296] = 8'b11110011;
mem1[3297] = 8'b11110011;
mem1[3298] = 8'b11110011;
mem1[3299] = 8'b11110011;
mem1[3300] = 8'b11110011;
mem1[3301] = 8'b11110011;
mem1[3302] = 8'b11110011;
mem1[3303] = 8'b11110011;
mem1[3304] = 8'b11110011;
mem1[3305] = 8'b11110011;
mem1[3306] = 8'b11110100;
mem1[3307] = 8'b11110100;
mem1[3308] = 8'b11110100;
mem1[3309] = 8'b11110100;
mem1[3310] = 8'b11110100;
mem1[3311] = 8'b11110100;
mem1[3312] = 8'b11110100;
mem1[3313] = 8'b11110100;
mem1[3314] = 8'b11110100;
mem1[3315] = 8'b11110100;
mem1[3316] = 8'b11110100;
mem1[3317] = 8'b11110100;
mem1[3318] = 8'b11110100;
mem1[3319] = 8'b11110100;
mem1[3320] = 8'b11110100;
mem1[3321] = 8'b11110100;
mem1[3322] = 8'b11110100;
mem1[3323] = 8'b11110100;
mem1[3324] = 8'b11110100;
mem1[3325] = 8'b11110100;
mem1[3326] = 8'b11110100;
mem1[3327] = 8'b11110100;
mem1[3328] = 8'b11110100;
mem1[3329] = 8'b11110101;
mem1[3330] = 8'b11110101;
mem1[3331] = 8'b11110101;
mem1[3332] = 8'b11110101;
mem1[3333] = 8'b11110101;
mem1[3334] = 8'b11110101;
mem1[3335] = 8'b11110101;
mem1[3336] = 8'b11110101;
mem1[3337] = 8'b11110101;
mem1[3338] = 8'b11110101;
mem1[3339] = 8'b11110101;
mem1[3340] = 8'b11110101;
mem1[3341] = 8'b11110101;
mem1[3342] = 8'b11110101;
mem1[3343] = 8'b11110101;
mem1[3344] = 8'b11110101;
mem1[3345] = 8'b11110101;
mem1[3346] = 8'b11110101;
mem1[3347] = 8'b11110101;
mem1[3348] = 8'b11110101;
mem1[3349] = 8'b11110101;
mem1[3350] = 8'b11110101;
mem1[3351] = 8'b11110101;
mem1[3352] = 8'b11110101;
mem1[3353] = 8'b11110110;
mem1[3354] = 8'b11110110;
mem1[3355] = 8'b11110110;
mem1[3356] = 8'b11110110;
mem1[3357] = 8'b11110110;
mem1[3358] = 8'b11110110;
mem1[3359] = 8'b11110110;
mem1[3360] = 8'b11110110;
mem1[3361] = 8'b11110110;
mem1[3362] = 8'b11110110;
mem1[3363] = 8'b11110110;
mem1[3364] = 8'b11110110;
mem1[3365] = 8'b11110110;
mem1[3366] = 8'b11110110;
mem1[3367] = 8'b11110110;
mem1[3368] = 8'b11110110;
mem1[3369] = 8'b11110110;
mem1[3370] = 8'b11110110;
mem1[3371] = 8'b11110110;
mem1[3372] = 8'b11110110;
mem1[3373] = 8'b11110110;
mem1[3374] = 8'b11110110;
mem1[3375] = 8'b11110110;
mem1[3376] = 8'b11110110;
mem1[3377] = 8'b11110110;
mem1[3378] = 8'b11110110;
mem1[3379] = 8'b11110111;
mem1[3380] = 8'b11110111;
mem1[3381] = 8'b11110111;
mem1[3382] = 8'b11110111;
mem1[3383] = 8'b11110111;
mem1[3384] = 8'b11110111;
mem1[3385] = 8'b11110111;
mem1[3386] = 8'b11110111;
mem1[3387] = 8'b11110111;
mem1[3388] = 8'b11110111;
mem1[3389] = 8'b11110111;
mem1[3390] = 8'b11110111;
mem1[3391] = 8'b11110111;
mem1[3392] = 8'b11110111;
mem1[3393] = 8'b11110111;
mem1[3394] = 8'b11110111;
mem1[3395] = 8'b11110111;
mem1[3396] = 8'b11110111;
mem1[3397] = 8'b11110111;
mem1[3398] = 8'b11110111;
mem1[3399] = 8'b11110111;
mem1[3400] = 8'b11110111;
mem1[3401] = 8'b11110111;
mem1[3402] = 8'b11110111;
mem1[3403] = 8'b11110111;
mem1[3404] = 8'b11110111;
mem1[3405] = 8'b11111000;
mem1[3406] = 8'b11111000;
mem1[3407] = 8'b11111000;
mem1[3408] = 8'b11111000;
mem1[3409] = 8'b11111000;
mem1[3410] = 8'b11111000;
mem1[3411] = 8'b11111000;
mem1[3412] = 8'b11111000;
mem1[3413] = 8'b11111000;
mem1[3414] = 8'b11111000;
mem1[3415] = 8'b11111000;
mem1[3416] = 8'b11111000;
mem1[3417] = 8'b11111000;
mem1[3418] = 8'b11111000;
mem1[3419] = 8'b11111000;
mem1[3420] = 8'b11111000;
mem1[3421] = 8'b11111000;
mem1[3422] = 8'b11111000;
mem1[3423] = 8'b11111000;
mem1[3424] = 8'b11111000;
mem1[3425] = 8'b11111000;
mem1[3426] = 8'b11111000;
mem1[3427] = 8'b11111000;
mem1[3428] = 8'b11111000;
mem1[3429] = 8'b11111000;
mem1[3430] = 8'b11111000;
mem1[3431] = 8'b11111000;
mem1[3432] = 8'b11111000;
mem1[3433] = 8'b11111000;
mem1[3434] = 8'b11111001;
mem1[3435] = 8'b11111001;
mem1[3436] = 8'b11111001;
mem1[3437] = 8'b11111001;
mem1[3438] = 8'b11111001;
mem1[3439] = 8'b11111001;
mem1[3440] = 8'b11111001;
mem1[3441] = 8'b11111001;
mem1[3442] = 8'b11111001;
mem1[3443] = 8'b11111001;
mem1[3444] = 8'b11111001;
mem1[3445] = 8'b11111001;
mem1[3446] = 8'b11111001;
mem1[3447] = 8'b11111001;
mem1[3448] = 8'b11111001;
mem1[3449] = 8'b11111001;
mem1[3450] = 8'b11111001;
mem1[3451] = 8'b11111001;
mem1[3452] = 8'b11111001;
mem1[3453] = 8'b11111001;
mem1[3454] = 8'b11111001;
mem1[3455] = 8'b11111001;
mem1[3456] = 8'b11111001;
mem1[3457] = 8'b11111001;
mem1[3458] = 8'b11111001;
mem1[3459] = 8'b11111001;
mem1[3460] = 8'b11111001;
mem1[3461] = 8'b11111001;
mem1[3462] = 8'b11111001;
mem1[3463] = 8'b11111001;
mem1[3464] = 8'b11111010;
mem1[3465] = 8'b11111010;
mem1[3466] = 8'b11111010;
mem1[3467] = 8'b11111010;
mem1[3468] = 8'b11111010;
mem1[3469] = 8'b11111010;
mem1[3470] = 8'b11111010;
mem1[3471] = 8'b11111010;
mem1[3472] = 8'b11111010;
mem1[3473] = 8'b11111010;
mem1[3474] = 8'b11111010;
mem1[3475] = 8'b11111010;
mem1[3476] = 8'b11111010;
mem1[3477] = 8'b11111010;
mem1[3478] = 8'b11111010;
mem1[3479] = 8'b11111010;
mem1[3480] = 8'b11111010;
mem1[3481] = 8'b11111010;
mem1[3482] = 8'b11111010;
mem1[3483] = 8'b11111010;
mem1[3484] = 8'b11111010;
mem1[3485] = 8'b11111010;
mem1[3486] = 8'b11111010;
mem1[3487] = 8'b11111010;
mem1[3488] = 8'b11111010;
mem1[3489] = 8'b11111010;
mem1[3490] = 8'b11111010;
mem1[3491] = 8'b11111010;
mem1[3492] = 8'b11111010;
mem1[3493] = 8'b11111010;
mem1[3494] = 8'b11111010;
mem1[3495] = 8'b11111010;
mem1[3496] = 8'b11111010;
mem1[3497] = 8'b11111011;
mem1[3498] = 8'b11111011;
mem1[3499] = 8'b11111011;
mem1[3500] = 8'b11111011;
mem1[3501] = 8'b11111011;
mem1[3502] = 8'b11111011;
mem1[3503] = 8'b11111011;
mem1[3504] = 8'b11111011;
mem1[3505] = 8'b11111011;
mem1[3506] = 8'b11111011;
mem1[3507] = 8'b11111011;
mem1[3508] = 8'b11111011;
mem1[3509] = 8'b11111011;
mem1[3510] = 8'b11111011;
mem1[3511] = 8'b11111011;
mem1[3512] = 8'b11111011;
mem1[3513] = 8'b11111011;
mem1[3514] = 8'b11111011;
mem1[3515] = 8'b11111011;
mem1[3516] = 8'b11111011;
mem1[3517] = 8'b11111011;
mem1[3518] = 8'b11111011;
mem1[3519] = 8'b11111011;
mem1[3520] = 8'b11111011;
mem1[3521] = 8'b11111011;
mem1[3522] = 8'b11111011;
mem1[3523] = 8'b11111011;
mem1[3524] = 8'b11111011;
mem1[3525] = 8'b11111011;
mem1[3526] = 8'b11111011;
mem1[3527] = 8'b11111011;
mem1[3528] = 8'b11111011;
mem1[3529] = 8'b11111011;
mem1[3530] = 8'b11111011;
mem1[3531] = 8'b11111011;
mem1[3532] = 8'b11111011;
mem1[3533] = 8'b11111100;
mem1[3534] = 8'b11111100;
mem1[3535] = 8'b11111100;
mem1[3536] = 8'b11111100;
mem1[3537] = 8'b11111100;
mem1[3538] = 8'b11111100;
mem1[3539] = 8'b11111100;
mem1[3540] = 8'b11111100;
mem1[3541] = 8'b11111100;
mem1[3542] = 8'b11111100;
mem1[3543] = 8'b11111100;
mem1[3544] = 8'b11111100;
mem1[3545] = 8'b11111100;
mem1[3546] = 8'b11111100;
mem1[3547] = 8'b11111100;
mem1[3548] = 8'b11111100;
mem1[3549] = 8'b11111100;
mem1[3550] = 8'b11111100;
mem1[3551] = 8'b11111100;
mem1[3552] = 8'b11111100;
mem1[3553] = 8'b11111100;
mem1[3554] = 8'b11111100;
mem1[3555] = 8'b11111100;
mem1[3556] = 8'b11111100;
mem1[3557] = 8'b11111100;
mem1[3558] = 8'b11111100;
mem1[3559] = 8'b11111100;
mem1[3560] = 8'b11111100;
mem1[3561] = 8'b11111100;
mem1[3562] = 8'b11111100;
mem1[3563] = 8'b11111100;
mem1[3564] = 8'b11111100;
mem1[3565] = 8'b11111100;
mem1[3566] = 8'b11111100;
mem1[3567] = 8'b11111100;
mem1[3568] = 8'b11111100;
mem1[3569] = 8'b11111100;
mem1[3570] = 8'b11111100;
mem1[3571] = 8'b11111100;
mem1[3572] = 8'b11111100;
mem1[3573] = 8'b11111100;
mem1[3574] = 8'b11111100;
mem1[3575] = 8'b11111101;
mem1[3576] = 8'b11111101;
mem1[3577] = 8'b11111101;
mem1[3578] = 8'b11111101;
mem1[3579] = 8'b11111101;
mem1[3580] = 8'b11111101;
mem1[3581] = 8'b11111101;
mem1[3582] = 8'b11111101;
mem1[3583] = 8'b11111101;
mem1[3584] = 8'b11111101;
mem1[3585] = 8'b11111101;
mem1[3586] = 8'b11111101;
mem1[3587] = 8'b11111101;
mem1[3588] = 8'b11111101;
mem1[3589] = 8'b11111101;
mem1[3590] = 8'b11111101;
mem1[3591] = 8'b11111101;
mem1[3592] = 8'b11111101;
mem1[3593] = 8'b11111101;
mem1[3594] = 8'b11111101;
mem1[3595] = 8'b11111101;
mem1[3596] = 8'b11111101;
mem1[3597] = 8'b11111101;
mem1[3598] = 8'b11111101;
mem1[3599] = 8'b11111101;
mem1[3600] = 8'b11111101;
mem1[3601] = 8'b11111101;
mem1[3602] = 8'b11111101;
mem1[3603] = 8'b11111101;
mem1[3604] = 8'b11111101;
mem1[3605] = 8'b11111101;
mem1[3606] = 8'b11111101;
mem1[3607] = 8'b11111101;
mem1[3608] = 8'b11111101;
mem1[3609] = 8'b11111101;
mem1[3610] = 8'b11111101;
mem1[3611] = 8'b11111101;
mem1[3612] = 8'b11111101;
mem1[3613] = 8'b11111101;
mem1[3614] = 8'b11111101;
mem1[3615] = 8'b11111101;
mem1[3616] = 8'b11111101;
mem1[3617] = 8'b11111101;
mem1[3618] = 8'b11111101;
mem1[3619] = 8'b11111101;
mem1[3620] = 8'b11111101;
mem1[3621] = 8'b11111101;
mem1[3622] = 8'b11111101;
mem1[3623] = 8'b11111110;
mem1[3624] = 8'b11111110;
mem1[3625] = 8'b11111110;
mem1[3626] = 8'b11111110;
mem1[3627] = 8'b11111110;
mem1[3628] = 8'b11111110;
mem1[3629] = 8'b11111110;
mem1[3630] = 8'b11111110;
mem1[3631] = 8'b11111110;
mem1[3632] = 8'b11111110;
mem1[3633] = 8'b11111110;
mem1[3634] = 8'b11111110;
mem1[3635] = 8'b11111110;
mem1[3636] = 8'b11111110;
mem1[3637] = 8'b11111110;
mem1[3638] = 8'b11111110;
mem1[3639] = 8'b11111110;
mem1[3640] = 8'b11111110;
mem1[3641] = 8'b11111110;
mem1[3642] = 8'b11111110;
mem1[3643] = 8'b11111110;
mem1[3644] = 8'b11111110;
mem1[3645] = 8'b11111110;
mem1[3646] = 8'b11111110;
mem1[3647] = 8'b11111110;
mem1[3648] = 8'b11111110;
mem1[3649] = 8'b11111110;
mem1[3650] = 8'b11111110;
mem1[3651] = 8'b11111110;
mem1[3652] = 8'b11111110;
mem1[3653] = 8'b11111110;
mem1[3654] = 8'b11111110;
mem1[3655] = 8'b11111110;
mem1[3656] = 8'b11111110;
mem1[3657] = 8'b11111110;
mem1[3658] = 8'b11111110;
mem1[3659] = 8'b11111110;
mem1[3660] = 8'b11111110;
mem1[3661] = 8'b11111110;
mem1[3662] = 8'b11111110;
mem1[3663] = 8'b11111110;
mem1[3664] = 8'b11111110;
mem1[3665] = 8'b11111110;
mem1[3666] = 8'b11111110;
mem1[3667] = 8'b11111110;
mem1[3668] = 8'b11111110;
mem1[3669] = 8'b11111110;
mem1[3670] = 8'b11111110;
mem1[3671] = 8'b11111110;
mem1[3672] = 8'b11111110;
mem1[3673] = 8'b11111110;
mem1[3674] = 8'b11111110;
mem1[3675] = 8'b11111110;
mem1[3676] = 8'b11111110;
mem1[3677] = 8'b11111110;
mem1[3678] = 8'b11111110;
mem1[3679] = 8'b11111110;
mem1[3680] = 8'b11111110;
mem1[3681] = 8'b11111110;
mem1[3682] = 8'b11111110;
mem1[3683] = 8'b11111110;
mem1[3684] = 8'b11111110;
mem1[3685] = 8'b11111110;
mem1[3686] = 8'b11111110;
mem1[3687] = 8'b11111111;
mem1[3688] = 8'b11111111;
mem1[3689] = 8'b11111111;
mem1[3690] = 8'b11111111;
mem1[3691] = 8'b11111111;
mem1[3692] = 8'b11111111;
mem1[3693] = 8'b11111111;
mem1[3694] = 8'b11111111;
mem1[3695] = 8'b11111111;
mem1[3696] = 8'b11111111;
mem1[3697] = 8'b11111111;
mem1[3698] = 8'b11111111;
mem1[3699] = 8'b11111111;
mem1[3700] = 8'b11111111;
mem1[3701] = 8'b11111111;
mem1[3702] = 8'b11111111;
mem1[3703] = 8'b11111111;
mem1[3704] = 8'b11111111;
mem1[3705] = 8'b11111111;
mem1[3706] = 8'b11111111;
mem1[3707] = 8'b11111111;
mem1[3708] = 8'b11111111;
mem1[3709] = 8'b11111111;
mem1[3710] = 8'b11111111;
mem1[3711] = 8'b11111111;
mem1[3712] = 8'b11111111;
mem1[3713] = 8'b11111111;
mem1[3714] = 8'b11111111;
mem1[3715] = 8'b11111111;
mem1[3716] = 8'b11111111;
mem1[3717] = 8'b11111111;
mem1[3718] = 8'b11111111;
mem1[3719] = 8'b11111111;
mem1[3720] = 8'b11111111;
mem1[3721] = 8'b11111111;
mem1[3722] = 8'b11111111;
mem1[3723] = 8'b11111111;
mem1[3724] = 8'b11111111;
mem1[3725] = 8'b11111111;
mem1[3726] = 8'b11111111;
mem1[3727] = 8'b11111111;
mem1[3728] = 8'b11111111;
mem1[3729] = 8'b11111111;
mem1[3730] = 8'b11111111;
mem1[3731] = 8'b11111111;
mem1[3732] = 8'b11111111;
mem1[3733] = 8'b11111111;
mem1[3734] = 8'b11111111;
mem1[3735] = 8'b11111111;
mem1[3736] = 8'b11111111;
mem1[3737] = 8'b11111111;
mem1[3738] = 8'b11111111;
mem1[3739] = 8'b11111111;
mem1[3740] = 8'b11111111;
mem1[3741] = 8'b11111111;
mem1[3742] = 8'b11111111;
mem1[3743] = 8'b11111111;
mem1[3744] = 8'b11111111;
mem1[3745] = 8'b11111111;
mem1[3746] = 8'b11111111;
mem1[3747] = 8'b11111111;
mem1[3748] = 8'b11111111;
mem1[3749] = 8'b11111111;
mem1[3750] = 8'b11111111;
mem1[3751] = 8'b11111111;
mem1[3752] = 8'b11111111;
mem1[3753] = 8'b11111111;
mem1[3754] = 8'b11111111;
mem1[3755] = 8'b11111111;
mem1[3756] = 8'b11111111;
mem1[3757] = 8'b11111111;
mem1[3758] = 8'b11111111;
mem1[3759] = 8'b11111111;
mem1[3760] = 8'b11111111;
mem1[3761] = 8'b11111111;
mem1[3762] = 8'b11111111;
mem1[3763] = 8'b11111111;
mem1[3764] = 8'b11111111;
mem1[3765] = 8'b11111111;
mem1[3766] = 8'b11111111;
mem1[3767] = 8'b11111111;
mem1[3768] = 8'b11111111;
mem1[3769] = 8'b11111111;
mem1[3770] = 8'b11111111;
mem1[3771] = 8'b11111111;
mem1[3772] = 8'b11111111;
mem1[3773] = 8'b11111111;
mem1[3774] = 8'b11111111;
mem1[3775] = 8'b11111111;
mem1[3776] = 8'b11111111;
mem1[3777] = 8'b11111111;
mem1[3778] = 8'b11111111;
mem1[3779] = 8'b11111111;
mem1[3780] = 8'b11111111;
mem1[3781] = 8'b11111111;
mem1[3782] = 8'b11111111;
mem1[3783] = 8'b11111111;
mem1[3784] = 8'b11111111;
mem1[3785] = 8'b11111111;
mem1[3786] = 8'b11111111;
mem1[3787] = 8'b11111111;
mem1[3788] = 8'b11111111;
mem1[3789] = 8'b11111111;
mem1[3790] = 8'b11111111;
mem1[3791] = 8'b11111111;
mem1[3792] = 8'b11111111;
mem1[3793] = 8'b11111111;
mem1[3794] = 8'b11111111;
mem1[3795] = 8'b11111111;
mem1[3796] = 8'b11111111;
mem1[3797] = 8'b11111111;
mem1[3798] = 8'b11111111;
mem1[3799] = 8'b11111111;
mem1[3800] = 8'b11111111;
mem1[3801] = 8'b11111111;
mem1[3802] = 8'b11111111;
mem1[3803] = 8'b11111111;
mem1[3804] = 8'b11111111;
mem1[3805] = 8'b11111111;
mem1[3806] = 8'b11111111;
mem1[3807] = 8'b11111111;
mem1[3808] = 8'b11111111;
mem1[3809] = 8'b11111111;
mem1[3810] = 8'b11111111;
mem1[3811] = 8'b11111111;
mem1[3812] = 8'b11111111;
mem1[3813] = 8'b11111111;
mem1[3814] = 8'b11111111;
mem1[3815] = 8'b11111111;
mem1[3816] = 8'b11111111;
mem1[3817] = 8'b11111111;
mem1[3818] = 8'b11111111;
mem1[3819] = 8'b11111111;
mem1[3820] = 8'b11111111;
mem1[3821] = 8'b11111111;
mem1[3822] = 8'b11111111;
mem1[3823] = 8'b11111111;
mem1[3824] = 8'b11111111;
mem1[3825] = 8'b11111111;
mem1[3826] = 8'b11111111;
mem1[3827] = 8'b11111111;
mem1[3828] = 8'b11111111;
mem1[3829] = 8'b11111111;
mem1[3830] = 8'b11111111;
mem1[3831] = 8'b11111111;
mem1[3832] = 8'b11111111;
mem1[3833] = 8'b11111111;
mem1[3834] = 8'b11111111;
mem1[3835] = 8'b11111111;
mem1[3836] = 8'b11111111;
mem1[3837] = 8'b11111111;
mem1[3838] = 8'b11111111;
mem1[3839] = 8'b11111111;
end

always @(posedge clk1) begin
	output_data_1 = mem1[selector1];
end

endmodule